`include "Parameter.v"
module Adder_tree 
(
   input   [`NBIT*`NDATA-1:0]    i_data,
   input   [`NDATA-1:0]    i_sign,
   output  [`NRESULT:0]          o_result
);

wire stage_0 [`NBIT-1:0][`NDATA*2:0];
genvar i, j;

generate
for (i=0; i<`NDATA; i=i+1) begin: i_loop_i_data
    for (j=0; j<`NBIT; j=j+1) begin: j_loop_i_data
       assign stage_0[j][i] = i_data[j+i*`NBIT];
    end;
end
endgenerate
generate
for (i=`NDATA; i<`NDATA*2; i=i+1) begin: i_loop_i_sign
    assign stage_0[0][i] = i_sign[i-`NDATA];
end
endgenerate


wire stage_1 [`NBIT+1:0][`NDATA*2:0];
FA FA_1_0 ( .a(stage_0[0][0]), .b(stage_0[0][1]), .cin(stage_0[0][2]), .cout(stage_1[1][0]), .s(stage_1[0][0]) );
FA FA_1_1 ( .a(stage_0[0][3]), .b(stage_0[0][4]), .cin(stage_0[0][5]), .cout(stage_1[1][1]), .s(stage_1[0][1]) );
FA FA_1_2 ( .a(stage_0[0][6]), .b(stage_0[0][7]), .cin(stage_0[0][8]), .cout(stage_1[1][2]), .s(stage_1[0][2]) );
FA FA_1_3 ( .a(stage_0[0][9]), .b(stage_0[0][10]), .cin(stage_0[0][11]), .cout(stage_1[1][3]), .s(stage_1[0][3]) );
FA FA_1_4 ( .a(stage_0[0][12]), .b(stage_0[0][13]), .cin(stage_0[0][14]), .cout(stage_1[1][4]), .s(stage_1[0][4]) );
FA FA_1_5 ( .a(stage_0[0][15]), .b(stage_0[0][16]), .cin(stage_0[0][17]), .cout(stage_1[1][5]), .s(stage_1[0][5]) );
FA FA_1_6 ( .a(stage_0[0][18]), .b(stage_0[0][19]), .cin(stage_0[0][20]), .cout(stage_1[1][6]), .s(stage_1[0][6]) );
FA FA_1_7 ( .a(stage_0[0][21]), .b(stage_0[0][22]), .cin(stage_0[0][23]), .cout(stage_1[1][7]), .s(stage_1[0][7]) );
FA FA_1_8 ( .a(stage_0[0][24]), .b(stage_0[0][25]), .cin(stage_0[0][26]), .cout(stage_1[1][8]), .s(stage_1[0][8]) );
FA FA_1_9 ( .a(stage_0[0][27]), .b(stage_0[0][28]), .cin(stage_0[0][29]), .cout(stage_1[1][9]), .s(stage_1[0][9]) );
FA FA_1_10 ( .a(stage_0[0][30]), .b(stage_0[0][31]), .cin(stage_0[0][32]), .cout(stage_1[1][10]), .s(stage_1[0][10]) );
FA FA_1_11 ( .a(stage_0[0][33]), .b(stage_0[0][34]), .cin(stage_0[0][35]), .cout(stage_1[1][11]), .s(stage_1[0][11]) );
FA FA_1_12 ( .a(stage_0[0][36]), .b(stage_0[0][37]), .cin(stage_0[0][38]), .cout(stage_1[1][12]), .s(stage_1[0][12]) );
FA FA_1_13 ( .a(stage_0[0][39]), .b(stage_0[0][40]), .cin(stage_0[0][41]), .cout(stage_1[1][13]), .s(stage_1[0][13]) );
FA FA_1_14 ( .a(stage_0[0][42]), .b(stage_0[0][43]), .cin(stage_0[0][44]), .cout(stage_1[1][14]), .s(stage_1[0][14]) );
FA FA_1_15 ( .a(stage_0[0][45]), .b(stage_0[0][46]), .cin(stage_0[0][47]), .cout(stage_1[1][15]), .s(stage_1[0][15]) );
FA FA_1_16 ( .a(stage_0[0][48]), .b(stage_0[0][49]), .cin(stage_0[0][50]), .cout(stage_1[1][16]), .s(stage_1[0][16]) );
FA FA_1_17 ( .a(stage_0[0][51]), .b(stage_0[0][52]), .cin(stage_0[0][53]), .cout(stage_1[1][17]), .s(stage_1[0][17]) );
FA FA_1_18 ( .a(stage_0[0][54]), .b(stage_0[0][55]), .cin(stage_0[0][56]), .cout(stage_1[1][18]), .s(stage_1[0][18]) );
FA FA_1_19 ( .a(stage_0[0][57]), .b(stage_0[0][58]), .cin(stage_0[0][59]), .cout(stage_1[1][19]), .s(stage_1[0][19]) );
FA FA_1_20 ( .a(stage_0[0][60]), .b(stage_0[0][61]), .cin(stage_0[0][62]), .cout(stage_1[1][20]), .s(stage_1[0][20]) );
FA FA_1_21 ( .a(stage_0[0][63]), .b(stage_0[0][64]), .cin(stage_0[0][65]), .cout(stage_1[1][21]), .s(stage_1[0][21]) );
FA FA_1_22 ( .a(stage_0[0][66]), .b(stage_0[0][67]), .cin(stage_0[0][68]), .cout(stage_1[1][22]), .s(stage_1[0][22]) );
FA FA_1_23 ( .a(stage_0[0][69]), .b(stage_0[0][70]), .cin(stage_0[0][71]), .cout(stage_1[1][23]), .s(stage_1[0][23]) );
FA FA_1_24 ( .a(stage_0[0][72]), .b(stage_0[0][73]), .cin(stage_0[0][74]), .cout(stage_1[1][24]), .s(stage_1[0][24]) );
FA FA_1_25 ( .a(stage_0[0][75]), .b(stage_0[0][76]), .cin(stage_0[0][77]), .cout(stage_1[1][25]), .s(stage_1[0][25]) );
FA FA_1_26 ( .a(stage_0[0][78]), .b(stage_0[0][79]), .cin(stage_0[0][80]), .cout(stage_1[1][26]), .s(stage_1[0][26]) );
FA FA_1_27 ( .a(stage_0[0][81]), .b(stage_0[0][82]), .cin(stage_0[0][83]), .cout(stage_1[1][27]), .s(stage_1[0][27]) );
FA FA_1_28 ( .a(stage_0[0][84]), .b(stage_0[0][85]), .cin(stage_0[0][86]), .cout(stage_1[1][28]), .s(stage_1[0][28]) );
FA FA_1_29 ( .a(stage_0[0][87]), .b(stage_0[0][88]), .cin(stage_0[0][89]), .cout(stage_1[1][29]), .s(stage_1[0][29]) );
FA FA_1_30 ( .a(stage_0[0][90]), .b(stage_0[0][91]), .cin(stage_0[0][92]), .cout(stage_1[1][30]), .s(stage_1[0][30]) );
FA FA_1_31 ( .a(stage_0[0][93]), .b(stage_0[0][94]), .cin(stage_0[0][95]), .cout(stage_1[1][31]), .s(stage_1[0][31]) );
FA FA_1_32 ( .a(stage_0[0][96]), .b(stage_0[0][97]), .cin(stage_0[0][98]), .cout(stage_1[1][32]), .s(stage_1[0][32]) );
FA FA_1_33 ( .a(stage_0[0][99]), .b(stage_0[0][100]), .cin(stage_0[0][101]), .cout(stage_1[1][33]), .s(stage_1[0][33]) );
FA FA_1_34 ( .a(stage_0[0][102]), .b(stage_0[0][103]), .cin(stage_0[0][104]), .cout(stage_1[1][34]), .s(stage_1[0][34]) );
FA FA_1_35 ( .a(stage_0[0][105]), .b(stage_0[0][106]), .cin(stage_0[0][107]), .cout(stage_1[1][35]), .s(stage_1[0][35]) );
FA FA_1_36 ( .a(stage_0[0][108]), .b(stage_0[0][109]), .cin(stage_0[0][110]), .cout(stage_1[1][36]), .s(stage_1[0][36]) );
FA FA_1_37 ( .a(stage_0[0][111]), .b(stage_0[0][112]), .cin(stage_0[0][113]), .cout(stage_1[1][37]), .s(stage_1[0][37]) );
FA FA_1_38 ( .a(stage_0[0][114]), .b(stage_0[0][115]), .cin(stage_0[0][116]), .cout(stage_1[1][38]), .s(stage_1[0][38]) );
FA FA_1_39 ( .a(stage_0[0][117]), .b(stage_0[0][118]), .cin(stage_0[0][119]), .cout(stage_1[1][39]), .s(stage_1[0][39]) );
FA FA_1_40 ( .a(stage_0[0][120]), .b(stage_0[0][121]), .cin(stage_0[0][122]), .cout(stage_1[1][40]), .s(stage_1[0][40]) );
FA FA_1_41 ( .a(stage_0[0][123]), .b(stage_0[0][124]), .cin(stage_0[0][125]), .cout(stage_1[1][41]), .s(stage_1[0][41]) );
HA HA_1_0 ( .a(stage_0[0][126]), .b(stage_0[0][127]), .cout(stage_1[1][42]), .s(stage_1[0][42]) );
FA FA_1_42 ( .a(stage_0[1][0]), .b(stage_0[1][1]), .cin(stage_0[1][2]), .cout(stage_1[2][0]), .s(stage_1[1][43]) );
FA FA_1_43 ( .a(stage_0[1][3]), .b(stage_0[1][4]), .cin(stage_0[1][5]), .cout(stage_1[2][1]), .s(stage_1[1][44]) );
FA FA_1_44 ( .a(stage_0[1][6]), .b(stage_0[1][7]), .cin(stage_0[1][8]), .cout(stage_1[2][2]), .s(stage_1[1][45]) );
FA FA_1_45 ( .a(stage_0[1][9]), .b(stage_0[1][10]), .cin(stage_0[1][11]), .cout(stage_1[2][3]), .s(stage_1[1][46]) );
FA FA_1_46 ( .a(stage_0[1][12]), .b(stage_0[1][13]), .cin(stage_0[1][14]), .cout(stage_1[2][4]), .s(stage_1[1][47]) );
FA FA_1_47 ( .a(stage_0[1][15]), .b(stage_0[1][16]), .cin(stage_0[1][17]), .cout(stage_1[2][5]), .s(stage_1[1][48]) );
FA FA_1_48 ( .a(stage_0[1][18]), .b(stage_0[1][19]), .cin(stage_0[1][20]), .cout(stage_1[2][6]), .s(stage_1[1][49]) );
FA FA_1_49 ( .a(stage_0[1][21]), .b(stage_0[1][22]), .cin(stage_0[1][23]), .cout(stage_1[2][7]), .s(stage_1[1][50]) );
FA FA_1_50 ( .a(stage_0[1][24]), .b(stage_0[1][25]), .cin(stage_0[1][26]), .cout(stage_1[2][8]), .s(stage_1[1][51]) );
FA FA_1_51 ( .a(stage_0[1][27]), .b(stage_0[1][28]), .cin(stage_0[1][29]), .cout(stage_1[2][9]), .s(stage_1[1][52]) );
FA FA_1_52 ( .a(stage_0[1][30]), .b(stage_0[1][31]), .cin(stage_0[1][32]), .cout(stage_1[2][10]), .s(stage_1[1][53]) );
FA FA_1_53 ( .a(stage_0[1][33]), .b(stage_0[1][34]), .cin(stage_0[1][35]), .cout(stage_1[2][11]), .s(stage_1[1][54]) );
FA FA_1_54 ( .a(stage_0[1][36]), .b(stage_0[1][37]), .cin(stage_0[1][38]), .cout(stage_1[2][12]), .s(stage_1[1][55]) );
FA FA_1_55 ( .a(stage_0[1][39]), .b(stage_0[1][40]), .cin(stage_0[1][41]), .cout(stage_1[2][13]), .s(stage_1[1][56]) );
FA FA_1_56 ( .a(stage_0[1][42]), .b(stage_0[1][43]), .cin(stage_0[1][44]), .cout(stage_1[2][14]), .s(stage_1[1][57]) );
FA FA_1_57 ( .a(stage_0[1][45]), .b(stage_0[1][46]), .cin(stage_0[1][47]), .cout(stage_1[2][15]), .s(stage_1[1][58]) );
FA FA_1_58 ( .a(stage_0[1][48]), .b(stage_0[1][49]), .cin(stage_0[1][50]), .cout(stage_1[2][16]), .s(stage_1[1][59]) );
FA FA_1_59 ( .a(stage_0[1][51]), .b(stage_0[1][52]), .cin(stage_0[1][53]), .cout(stage_1[2][17]), .s(stage_1[1][60]) );
FA FA_1_60 ( .a(stage_0[1][54]), .b(stage_0[1][55]), .cin(stage_0[1][56]), .cout(stage_1[2][18]), .s(stage_1[1][61]) );
FA FA_1_61 ( .a(stage_0[1][57]), .b(stage_0[1][58]), .cin(stage_0[1][59]), .cout(stage_1[2][19]), .s(stage_1[1][62]) );
FA FA_1_62 ( .a(stage_0[1][60]), .b(stage_0[1][61]), .cin(stage_0[1][62]), .cout(stage_1[2][20]), .s(stage_1[1][63]) );
assign stage_1[1][64] = stage_0[1][63];
FA FA_1_63 ( .a(stage_0[2][0]), .b(stage_0[2][1]), .cin(stage_0[2][2]), .cout(stage_1[3][0]), .s(stage_1[2][21]) );
FA FA_1_64 ( .a(stage_0[2][3]), .b(stage_0[2][4]), .cin(stage_0[2][5]), .cout(stage_1[3][1]), .s(stage_1[2][22]) );
FA FA_1_65 ( .a(stage_0[2][6]), .b(stage_0[2][7]), .cin(stage_0[2][8]), .cout(stage_1[3][2]), .s(stage_1[2][23]) );
FA FA_1_66 ( .a(stage_0[2][9]), .b(stage_0[2][10]), .cin(stage_0[2][11]), .cout(stage_1[3][3]), .s(stage_1[2][24]) );
FA FA_1_67 ( .a(stage_0[2][12]), .b(stage_0[2][13]), .cin(stage_0[2][14]), .cout(stage_1[3][4]), .s(stage_1[2][25]) );
FA FA_1_68 ( .a(stage_0[2][15]), .b(stage_0[2][16]), .cin(stage_0[2][17]), .cout(stage_1[3][5]), .s(stage_1[2][26]) );
FA FA_1_69 ( .a(stage_0[2][18]), .b(stage_0[2][19]), .cin(stage_0[2][20]), .cout(stage_1[3][6]), .s(stage_1[2][27]) );
FA FA_1_70 ( .a(stage_0[2][21]), .b(stage_0[2][22]), .cin(stage_0[2][23]), .cout(stage_1[3][7]), .s(stage_1[2][28]) );
FA FA_1_71 ( .a(stage_0[2][24]), .b(stage_0[2][25]), .cin(stage_0[2][26]), .cout(stage_1[3][8]), .s(stage_1[2][29]) );
FA FA_1_72 ( .a(stage_0[2][27]), .b(stage_0[2][28]), .cin(stage_0[2][29]), .cout(stage_1[3][9]), .s(stage_1[2][30]) );
FA FA_1_73 ( .a(stage_0[2][30]), .b(stage_0[2][31]), .cin(stage_0[2][32]), .cout(stage_1[3][10]), .s(stage_1[2][31]) );
FA FA_1_74 ( .a(stage_0[2][33]), .b(stage_0[2][34]), .cin(stage_0[2][35]), .cout(stage_1[3][11]), .s(stage_1[2][32]) );
FA FA_1_75 ( .a(stage_0[2][36]), .b(stage_0[2][37]), .cin(stage_0[2][38]), .cout(stage_1[3][12]), .s(stage_1[2][33]) );
FA FA_1_76 ( .a(stage_0[2][39]), .b(stage_0[2][40]), .cin(stage_0[2][41]), .cout(stage_1[3][13]), .s(stage_1[2][34]) );
FA FA_1_77 ( .a(stage_0[2][42]), .b(stage_0[2][43]), .cin(stage_0[2][44]), .cout(stage_1[3][14]), .s(stage_1[2][35]) );
FA FA_1_78 ( .a(stage_0[2][45]), .b(stage_0[2][46]), .cin(stage_0[2][47]), .cout(stage_1[3][15]), .s(stage_1[2][36]) );
FA FA_1_79 ( .a(stage_0[2][48]), .b(stage_0[2][49]), .cin(stage_0[2][50]), .cout(stage_1[3][16]), .s(stage_1[2][37]) );
FA FA_1_80 ( .a(stage_0[2][51]), .b(stage_0[2][52]), .cin(stage_0[2][53]), .cout(stage_1[3][17]), .s(stage_1[2][38]) );
FA FA_1_81 ( .a(stage_0[2][54]), .b(stage_0[2][55]), .cin(stage_0[2][56]), .cout(stage_1[3][18]), .s(stage_1[2][39]) );
FA FA_1_82 ( .a(stage_0[2][57]), .b(stage_0[2][58]), .cin(stage_0[2][59]), .cout(stage_1[3][19]), .s(stage_1[2][40]) );
FA FA_1_83 ( .a(stage_0[2][60]), .b(stage_0[2][61]), .cin(stage_0[2][62]), .cout(stage_1[3][20]), .s(stage_1[2][41]) );
assign stage_1[2][42] = stage_0[2][63];
FA FA_1_84 ( .a(stage_0[3][0]), .b(stage_0[3][1]), .cin(stage_0[3][2]), .cout(stage_1[4][0]), .s(stage_1[3][21]) );
FA FA_1_85 ( .a(stage_0[3][3]), .b(stage_0[3][4]), .cin(stage_0[3][5]), .cout(stage_1[4][1]), .s(stage_1[3][22]) );
FA FA_1_86 ( .a(stage_0[3][6]), .b(stage_0[3][7]), .cin(stage_0[3][8]), .cout(stage_1[4][2]), .s(stage_1[3][23]) );
FA FA_1_87 ( .a(stage_0[3][9]), .b(stage_0[3][10]), .cin(stage_0[3][11]), .cout(stage_1[4][3]), .s(stage_1[3][24]) );
FA FA_1_88 ( .a(stage_0[3][12]), .b(stage_0[3][13]), .cin(stage_0[3][14]), .cout(stage_1[4][4]), .s(stage_1[3][25]) );
FA FA_1_89 ( .a(stage_0[3][15]), .b(stage_0[3][16]), .cin(stage_0[3][17]), .cout(stage_1[4][5]), .s(stage_1[3][26]) );
FA FA_1_90 ( .a(stage_0[3][18]), .b(stage_0[3][19]), .cin(stage_0[3][20]), .cout(stage_1[4][6]), .s(stage_1[3][27]) );
FA FA_1_91 ( .a(stage_0[3][21]), .b(stage_0[3][22]), .cin(stage_0[3][23]), .cout(stage_1[4][7]), .s(stage_1[3][28]) );
FA FA_1_92 ( .a(stage_0[3][24]), .b(stage_0[3][25]), .cin(stage_0[3][26]), .cout(stage_1[4][8]), .s(stage_1[3][29]) );
FA FA_1_93 ( .a(stage_0[3][27]), .b(stage_0[3][28]), .cin(stage_0[3][29]), .cout(stage_1[4][9]), .s(stage_1[3][30]) );
FA FA_1_94 ( .a(stage_0[3][30]), .b(stage_0[3][31]), .cin(stage_0[3][32]), .cout(stage_1[4][10]), .s(stage_1[3][31]) );
FA FA_1_95 ( .a(stage_0[3][33]), .b(stage_0[3][34]), .cin(stage_0[3][35]), .cout(stage_1[4][11]), .s(stage_1[3][32]) );
FA FA_1_96 ( .a(stage_0[3][36]), .b(stage_0[3][37]), .cin(stage_0[3][38]), .cout(stage_1[4][12]), .s(stage_1[3][33]) );
FA FA_1_97 ( .a(stage_0[3][39]), .b(stage_0[3][40]), .cin(stage_0[3][41]), .cout(stage_1[4][13]), .s(stage_1[3][34]) );
FA FA_1_98 ( .a(stage_0[3][42]), .b(stage_0[3][43]), .cin(stage_0[3][44]), .cout(stage_1[4][14]), .s(stage_1[3][35]) );
FA FA_1_99 ( .a(stage_0[3][45]), .b(stage_0[3][46]), .cin(stage_0[3][47]), .cout(stage_1[4][15]), .s(stage_1[3][36]) );
FA FA_1_100 ( .a(stage_0[3][48]), .b(stage_0[3][49]), .cin(stage_0[3][50]), .cout(stage_1[4][16]), .s(stage_1[3][37]) );
FA FA_1_101 ( .a(stage_0[3][51]), .b(stage_0[3][52]), .cin(stage_0[3][53]), .cout(stage_1[4][17]), .s(stage_1[3][38]) );
FA FA_1_102 ( .a(stage_0[3][54]), .b(stage_0[3][55]), .cin(stage_0[3][56]), .cout(stage_1[4][18]), .s(stage_1[3][39]) );
FA FA_1_103 ( .a(stage_0[3][57]), .b(stage_0[3][58]), .cin(stage_0[3][59]), .cout(stage_1[4][19]), .s(stage_1[3][40]) );
FA FA_1_104 ( .a(stage_0[3][60]), .b(stage_0[3][61]), .cin(stage_0[3][62]), .cout(stage_1[4][20]), .s(stage_1[3][41]) );
assign stage_1[3][42] = stage_0[3][63];
FA FA_1_105 ( .a(stage_0[4][0]), .b(stage_0[4][1]), .cin(stage_0[4][2]), .cout(stage_1[5][0]), .s(stage_1[4][21]) );
FA FA_1_106 ( .a(stage_0[4][3]), .b(stage_0[4][4]), .cin(stage_0[4][5]), .cout(stage_1[5][1]), .s(stage_1[4][22]) );
FA FA_1_107 ( .a(stage_0[4][6]), .b(stage_0[4][7]), .cin(stage_0[4][8]), .cout(stage_1[5][2]), .s(stage_1[4][23]) );
FA FA_1_108 ( .a(stage_0[4][9]), .b(stage_0[4][10]), .cin(stage_0[4][11]), .cout(stage_1[5][3]), .s(stage_1[4][24]) );
FA FA_1_109 ( .a(stage_0[4][12]), .b(stage_0[4][13]), .cin(stage_0[4][14]), .cout(stage_1[5][4]), .s(stage_1[4][25]) );
FA FA_1_110 ( .a(stage_0[4][15]), .b(stage_0[4][16]), .cin(stage_0[4][17]), .cout(stage_1[5][5]), .s(stage_1[4][26]) );
FA FA_1_111 ( .a(stage_0[4][18]), .b(stage_0[4][19]), .cin(stage_0[4][20]), .cout(stage_1[5][6]), .s(stage_1[4][27]) );
FA FA_1_112 ( .a(stage_0[4][21]), .b(stage_0[4][22]), .cin(stage_0[4][23]), .cout(stage_1[5][7]), .s(stage_1[4][28]) );
FA FA_1_113 ( .a(stage_0[4][24]), .b(stage_0[4][25]), .cin(stage_0[4][26]), .cout(stage_1[5][8]), .s(stage_1[4][29]) );
FA FA_1_114 ( .a(stage_0[4][27]), .b(stage_0[4][28]), .cin(stage_0[4][29]), .cout(stage_1[5][9]), .s(stage_1[4][30]) );
FA FA_1_115 ( .a(stage_0[4][30]), .b(stage_0[4][31]), .cin(stage_0[4][32]), .cout(stage_1[5][10]), .s(stage_1[4][31]) );
FA FA_1_116 ( .a(stage_0[4][33]), .b(stage_0[4][34]), .cin(stage_0[4][35]), .cout(stage_1[5][11]), .s(stage_1[4][32]) );
FA FA_1_117 ( .a(stage_0[4][36]), .b(stage_0[4][37]), .cin(stage_0[4][38]), .cout(stage_1[5][12]), .s(stage_1[4][33]) );
FA FA_1_118 ( .a(stage_0[4][39]), .b(stage_0[4][40]), .cin(stage_0[4][41]), .cout(stage_1[5][13]), .s(stage_1[4][34]) );
FA FA_1_119 ( .a(stage_0[4][42]), .b(stage_0[4][43]), .cin(stage_0[4][44]), .cout(stage_1[5][14]), .s(stage_1[4][35]) );
FA FA_1_120 ( .a(stage_0[4][45]), .b(stage_0[4][46]), .cin(stage_0[4][47]), .cout(stage_1[5][15]), .s(stage_1[4][36]) );
FA FA_1_121 ( .a(stage_0[4][48]), .b(stage_0[4][49]), .cin(stage_0[4][50]), .cout(stage_1[5][16]), .s(stage_1[4][37]) );
FA FA_1_122 ( .a(stage_0[4][51]), .b(stage_0[4][52]), .cin(stage_0[4][53]), .cout(stage_1[5][17]), .s(stage_1[4][38]) );
FA FA_1_123 ( .a(stage_0[4][54]), .b(stage_0[4][55]), .cin(stage_0[4][56]), .cout(stage_1[5][18]), .s(stage_1[4][39]) );
FA FA_1_124 ( .a(stage_0[4][57]), .b(stage_0[4][58]), .cin(stage_0[4][59]), .cout(stage_1[5][19]), .s(stage_1[4][40]) );
FA FA_1_125 ( .a(stage_0[4][60]), .b(stage_0[4][61]), .cin(stage_0[4][62]), .cout(stage_1[5][20]), .s(stage_1[4][41]) );
assign stage_1[4][42] = stage_0[4][63];
FA FA_1_126 ( .a(stage_0[5][0]), .b(stage_0[5][1]), .cin(stage_0[5][2]), .cout(stage_1[6][0]), .s(stage_1[5][21]) );
FA FA_1_127 ( .a(stage_0[5][3]), .b(stage_0[5][4]), .cin(stage_0[5][5]), .cout(stage_1[6][1]), .s(stage_1[5][22]) );
FA FA_1_128 ( .a(stage_0[5][6]), .b(stage_0[5][7]), .cin(stage_0[5][8]), .cout(stage_1[6][2]), .s(stage_1[5][23]) );
FA FA_1_129 ( .a(stage_0[5][9]), .b(stage_0[5][10]), .cin(stage_0[5][11]), .cout(stage_1[6][3]), .s(stage_1[5][24]) );
FA FA_1_130 ( .a(stage_0[5][12]), .b(stage_0[5][13]), .cin(stage_0[5][14]), .cout(stage_1[6][4]), .s(stage_1[5][25]) );
FA FA_1_131 ( .a(stage_0[5][15]), .b(stage_0[5][16]), .cin(stage_0[5][17]), .cout(stage_1[6][5]), .s(stage_1[5][26]) );
FA FA_1_132 ( .a(stage_0[5][18]), .b(stage_0[5][19]), .cin(stage_0[5][20]), .cout(stage_1[6][6]), .s(stage_1[5][27]) );
FA FA_1_133 ( .a(stage_0[5][21]), .b(stage_0[5][22]), .cin(stage_0[5][23]), .cout(stage_1[6][7]), .s(stage_1[5][28]) );
FA FA_1_134 ( .a(stage_0[5][24]), .b(stage_0[5][25]), .cin(stage_0[5][26]), .cout(stage_1[6][8]), .s(stage_1[5][29]) );
FA FA_1_135 ( .a(stage_0[5][27]), .b(stage_0[5][28]), .cin(stage_0[5][29]), .cout(stage_1[6][9]), .s(stage_1[5][30]) );
FA FA_1_136 ( .a(stage_0[5][30]), .b(stage_0[5][31]), .cin(stage_0[5][32]), .cout(stage_1[6][10]), .s(stage_1[5][31]) );
FA FA_1_137 ( .a(stage_0[5][33]), .b(stage_0[5][34]), .cin(stage_0[5][35]), .cout(stage_1[6][11]), .s(stage_1[5][32]) );
FA FA_1_138 ( .a(stage_0[5][36]), .b(stage_0[5][37]), .cin(stage_0[5][38]), .cout(stage_1[6][12]), .s(stage_1[5][33]) );
FA FA_1_139 ( .a(stage_0[5][39]), .b(stage_0[5][40]), .cin(stage_0[5][41]), .cout(stage_1[6][13]), .s(stage_1[5][34]) );
FA FA_1_140 ( .a(stage_0[5][42]), .b(stage_0[5][43]), .cin(stage_0[5][44]), .cout(stage_1[6][14]), .s(stage_1[5][35]) );
FA FA_1_141 ( .a(stage_0[5][45]), .b(stage_0[5][46]), .cin(stage_0[5][47]), .cout(stage_1[6][15]), .s(stage_1[5][36]) );
FA FA_1_142 ( .a(stage_0[5][48]), .b(stage_0[5][49]), .cin(stage_0[5][50]), .cout(stage_1[6][16]), .s(stage_1[5][37]) );
FA FA_1_143 ( .a(stage_0[5][51]), .b(stage_0[5][52]), .cin(stage_0[5][53]), .cout(stage_1[6][17]), .s(stage_1[5][38]) );
FA FA_1_144 ( .a(stage_0[5][54]), .b(stage_0[5][55]), .cin(stage_0[5][56]), .cout(stage_1[6][18]), .s(stage_1[5][39]) );
FA FA_1_145 ( .a(stage_0[5][57]), .b(stage_0[5][58]), .cin(stage_0[5][59]), .cout(stage_1[6][19]), .s(stage_1[5][40]) );
FA FA_1_146 ( .a(stage_0[5][60]), .b(stage_0[5][61]), .cin(stage_0[5][62]), .cout(stage_1[6][20]), .s(stage_1[5][41]) );
assign stage_1[5][42] = stage_0[5][63];
FA FA_1_147 ( .a(stage_0[6][0]), .b(stage_0[6][1]), .cin(stage_0[6][2]), .cout(stage_1[7][0]), .s(stage_1[6][21]) );
FA FA_1_148 ( .a(stage_0[6][3]), .b(stage_0[6][4]), .cin(stage_0[6][5]), .cout(stage_1[7][1]), .s(stage_1[6][22]) );
FA FA_1_149 ( .a(stage_0[6][6]), .b(stage_0[6][7]), .cin(stage_0[6][8]), .cout(stage_1[7][2]), .s(stage_1[6][23]) );
FA FA_1_150 ( .a(stage_0[6][9]), .b(stage_0[6][10]), .cin(stage_0[6][11]), .cout(stage_1[7][3]), .s(stage_1[6][24]) );
FA FA_1_151 ( .a(stage_0[6][12]), .b(stage_0[6][13]), .cin(stage_0[6][14]), .cout(stage_1[7][4]), .s(stage_1[6][25]) );
FA FA_1_152 ( .a(stage_0[6][15]), .b(stage_0[6][16]), .cin(stage_0[6][17]), .cout(stage_1[7][5]), .s(stage_1[6][26]) );
FA FA_1_153 ( .a(stage_0[6][18]), .b(stage_0[6][19]), .cin(stage_0[6][20]), .cout(stage_1[7][6]), .s(stage_1[6][27]) );
FA FA_1_154 ( .a(stage_0[6][21]), .b(stage_0[6][22]), .cin(stage_0[6][23]), .cout(stage_1[7][7]), .s(stage_1[6][28]) );
FA FA_1_155 ( .a(stage_0[6][24]), .b(stage_0[6][25]), .cin(stage_0[6][26]), .cout(stage_1[7][8]), .s(stage_1[6][29]) );
FA FA_1_156 ( .a(stage_0[6][27]), .b(stage_0[6][28]), .cin(stage_0[6][29]), .cout(stage_1[7][9]), .s(stage_1[6][30]) );
FA FA_1_157 ( .a(stage_0[6][30]), .b(stage_0[6][31]), .cin(stage_0[6][32]), .cout(stage_1[7][10]), .s(stage_1[6][31]) );
FA FA_1_158 ( .a(stage_0[6][33]), .b(stage_0[6][34]), .cin(stage_0[6][35]), .cout(stage_1[7][11]), .s(stage_1[6][32]) );
FA FA_1_159 ( .a(stage_0[6][36]), .b(stage_0[6][37]), .cin(stage_0[6][38]), .cout(stage_1[7][12]), .s(stage_1[6][33]) );
FA FA_1_160 ( .a(stage_0[6][39]), .b(stage_0[6][40]), .cin(stage_0[6][41]), .cout(stage_1[7][13]), .s(stage_1[6][34]) );
FA FA_1_161 ( .a(stage_0[6][42]), .b(stage_0[6][43]), .cin(stage_0[6][44]), .cout(stage_1[7][14]), .s(stage_1[6][35]) );
FA FA_1_162 ( .a(stage_0[6][45]), .b(stage_0[6][46]), .cin(stage_0[6][47]), .cout(stage_1[7][15]), .s(stage_1[6][36]) );
FA FA_1_163 ( .a(stage_0[6][48]), .b(stage_0[6][49]), .cin(stage_0[6][50]), .cout(stage_1[7][16]), .s(stage_1[6][37]) );
FA FA_1_164 ( .a(stage_0[6][51]), .b(stage_0[6][52]), .cin(stage_0[6][53]), .cout(stage_1[7][17]), .s(stage_1[6][38]) );
FA FA_1_165 ( .a(stage_0[6][54]), .b(stage_0[6][55]), .cin(stage_0[6][56]), .cout(stage_1[7][18]), .s(stage_1[6][39]) );
FA FA_1_166 ( .a(stage_0[6][57]), .b(stage_0[6][58]), .cin(stage_0[6][59]), .cout(stage_1[7][19]), .s(stage_1[6][40]) );
FA FA_1_167 ( .a(stage_0[6][60]), .b(stage_0[6][61]), .cin(stage_0[6][62]), .cout(stage_1[7][20]), .s(stage_1[6][41]) );
assign stage_1[6][42] = stage_0[6][63];
FA FA_1_168 ( .a(stage_0[7][0]), .b(stage_0[7][1]), .cin(stage_0[7][2]), .cout(stage_1[8][0]), .s(stage_1[7][21]) );
FA FA_1_169 ( .a(stage_0[7][3]), .b(stage_0[7][4]), .cin(stage_0[7][5]), .cout(stage_1[8][1]), .s(stage_1[7][22]) );
FA FA_1_170 ( .a(stage_0[7][6]), .b(stage_0[7][7]), .cin(stage_0[7][8]), .cout(stage_1[8][2]), .s(stage_1[7][23]) );
FA FA_1_171 ( .a(stage_0[7][9]), .b(stage_0[7][10]), .cin(stage_0[7][11]), .cout(stage_1[8][3]), .s(stage_1[7][24]) );
FA FA_1_172 ( .a(stage_0[7][12]), .b(stage_0[7][13]), .cin(stage_0[7][14]), .cout(stage_1[8][4]), .s(stage_1[7][25]) );
FA FA_1_173 ( .a(stage_0[7][15]), .b(stage_0[7][16]), .cin(stage_0[7][17]), .cout(stage_1[8][5]), .s(stage_1[7][26]) );
FA FA_1_174 ( .a(stage_0[7][18]), .b(stage_0[7][19]), .cin(stage_0[7][20]), .cout(stage_1[8][6]), .s(stage_1[7][27]) );
FA FA_1_175 ( .a(stage_0[7][21]), .b(stage_0[7][22]), .cin(stage_0[7][23]), .cout(stage_1[8][7]), .s(stage_1[7][28]) );
FA FA_1_176 ( .a(stage_0[7][24]), .b(stage_0[7][25]), .cin(stage_0[7][26]), .cout(stage_1[8][8]), .s(stage_1[7][29]) );
FA FA_1_177 ( .a(stage_0[7][27]), .b(stage_0[7][28]), .cin(stage_0[7][29]), .cout(stage_1[8][9]), .s(stage_1[7][30]) );
FA FA_1_178 ( .a(stage_0[7][30]), .b(stage_0[7][31]), .cin(stage_0[7][32]), .cout(stage_1[8][10]), .s(stage_1[7][31]) );
FA FA_1_179 ( .a(stage_0[7][33]), .b(stage_0[7][34]), .cin(stage_0[7][35]), .cout(stage_1[8][11]), .s(stage_1[7][32]) );
FA FA_1_180 ( .a(stage_0[7][36]), .b(stage_0[7][37]), .cin(stage_0[7][38]), .cout(stage_1[8][12]), .s(stage_1[7][33]) );
FA FA_1_181 ( .a(stage_0[7][39]), .b(stage_0[7][40]), .cin(stage_0[7][41]), .cout(stage_1[8][13]), .s(stage_1[7][34]) );
FA FA_1_182 ( .a(stage_0[7][42]), .b(stage_0[7][43]), .cin(stage_0[7][44]), .cout(stage_1[8][14]), .s(stage_1[7][35]) );
FA FA_1_183 ( .a(stage_0[7][45]), .b(stage_0[7][46]), .cin(stage_0[7][47]), .cout(stage_1[8][15]), .s(stage_1[7][36]) );
FA FA_1_184 ( .a(stage_0[7][48]), .b(stage_0[7][49]), .cin(stage_0[7][50]), .cout(stage_1[8][16]), .s(stage_1[7][37]) );
FA FA_1_185 ( .a(stage_0[7][51]), .b(stage_0[7][52]), .cin(stage_0[7][53]), .cout(stage_1[8][17]), .s(stage_1[7][38]) );
FA FA_1_186 ( .a(stage_0[7][54]), .b(stage_0[7][55]), .cin(stage_0[7][56]), .cout(stage_1[8][18]), .s(stage_1[7][39]) );
FA FA_1_187 ( .a(stage_0[7][57]), .b(stage_0[7][58]), .cin(stage_0[7][59]), .cout(stage_1[8][19]), .s(stage_1[7][40]) );
FA FA_1_188 ( .a(stage_0[7][60]), .b(stage_0[7][61]), .cin(stage_0[7][62]), .cout(stage_1[8][20]), .s(stage_1[7][41]) );
assign stage_1[7][42] = stage_0[7][63];
FA FA_1_189 ( .a(stage_0[8][0]), .b(stage_0[8][1]), .cin(stage_0[8][2]), .cout(stage_1[9][0]), .s(stage_1[8][21]) );
FA FA_1_190 ( .a(stage_0[8][3]), .b(stage_0[8][4]), .cin(stage_0[8][5]), .cout(stage_1[9][1]), .s(stage_1[8][22]) );
FA FA_1_191 ( .a(stage_0[8][6]), .b(stage_0[8][7]), .cin(stage_0[8][8]), .cout(stage_1[9][2]), .s(stage_1[8][23]) );
FA FA_1_192 ( .a(stage_0[8][9]), .b(stage_0[8][10]), .cin(stage_0[8][11]), .cout(stage_1[9][3]), .s(stage_1[8][24]) );
FA FA_1_193 ( .a(stage_0[8][12]), .b(stage_0[8][13]), .cin(stage_0[8][14]), .cout(stage_1[9][4]), .s(stage_1[8][25]) );
FA FA_1_194 ( .a(stage_0[8][15]), .b(stage_0[8][16]), .cin(stage_0[8][17]), .cout(stage_1[9][5]), .s(stage_1[8][26]) );
FA FA_1_195 ( .a(stage_0[8][18]), .b(stage_0[8][19]), .cin(stage_0[8][20]), .cout(stage_1[9][6]), .s(stage_1[8][27]) );
FA FA_1_196 ( .a(stage_0[8][21]), .b(stage_0[8][22]), .cin(stage_0[8][23]), .cout(stage_1[9][7]), .s(stage_1[8][28]) );
FA FA_1_197 ( .a(stage_0[8][24]), .b(stage_0[8][25]), .cin(stage_0[8][26]), .cout(stage_1[9][8]), .s(stage_1[8][29]) );
FA FA_1_198 ( .a(stage_0[8][27]), .b(stage_0[8][28]), .cin(stage_0[8][29]), .cout(stage_1[9][9]), .s(stage_1[8][30]) );
FA FA_1_199 ( .a(stage_0[8][30]), .b(stage_0[8][31]), .cin(stage_0[8][32]), .cout(stage_1[9][10]), .s(stage_1[8][31]) );
FA FA_1_200 ( .a(stage_0[8][33]), .b(stage_0[8][34]), .cin(stage_0[8][35]), .cout(stage_1[9][11]), .s(stage_1[8][32]) );
FA FA_1_201 ( .a(stage_0[8][36]), .b(stage_0[8][37]), .cin(stage_0[8][38]), .cout(stage_1[9][12]), .s(stage_1[8][33]) );
FA FA_1_202 ( .a(stage_0[8][39]), .b(stage_0[8][40]), .cin(stage_0[8][41]), .cout(stage_1[9][13]), .s(stage_1[8][34]) );
FA FA_1_203 ( .a(stage_0[8][42]), .b(stage_0[8][43]), .cin(stage_0[8][44]), .cout(stage_1[9][14]), .s(stage_1[8][35]) );
FA FA_1_204 ( .a(stage_0[8][45]), .b(stage_0[8][46]), .cin(stage_0[8][47]), .cout(stage_1[9][15]), .s(stage_1[8][36]) );
FA FA_1_205 ( .a(stage_0[8][48]), .b(stage_0[8][49]), .cin(stage_0[8][50]), .cout(stage_1[9][16]), .s(stage_1[8][37]) );
FA FA_1_206 ( .a(stage_0[8][51]), .b(stage_0[8][52]), .cin(stage_0[8][53]), .cout(stage_1[9][17]), .s(stage_1[8][38]) );
FA FA_1_207 ( .a(stage_0[8][54]), .b(stage_0[8][55]), .cin(stage_0[8][56]), .cout(stage_1[9][18]), .s(stage_1[8][39]) );
FA FA_1_208 ( .a(stage_0[8][57]), .b(stage_0[8][58]), .cin(stage_0[8][59]), .cout(stage_1[9][19]), .s(stage_1[8][40]) );
FA FA_1_209 ( .a(stage_0[8][60]), .b(stage_0[8][61]), .cin(stage_0[8][62]), .cout(stage_1[9][20]), .s(stage_1[8][41]) );
assign stage_1[8][42] = stage_0[8][63];
FA FA_1_210 ( .a(stage_0[9][0]), .b(stage_0[9][1]), .cin(stage_0[9][2]), .cout(stage_1[10][0]), .s(stage_1[9][21]) );
FA FA_1_211 ( .a(stage_0[9][3]), .b(stage_0[9][4]), .cin(stage_0[9][5]), .cout(stage_1[10][1]), .s(stage_1[9][22]) );
FA FA_1_212 ( .a(stage_0[9][6]), .b(stage_0[9][7]), .cin(stage_0[9][8]), .cout(stage_1[10][2]), .s(stage_1[9][23]) );
FA FA_1_213 ( .a(stage_0[9][9]), .b(stage_0[9][10]), .cin(stage_0[9][11]), .cout(stage_1[10][3]), .s(stage_1[9][24]) );
FA FA_1_214 ( .a(stage_0[9][12]), .b(stage_0[9][13]), .cin(stage_0[9][14]), .cout(stage_1[10][4]), .s(stage_1[9][25]) );
FA FA_1_215 ( .a(stage_0[9][15]), .b(stage_0[9][16]), .cin(stage_0[9][17]), .cout(stage_1[10][5]), .s(stage_1[9][26]) );
FA FA_1_216 ( .a(stage_0[9][18]), .b(stage_0[9][19]), .cin(stage_0[9][20]), .cout(stage_1[10][6]), .s(stage_1[9][27]) );
FA FA_1_217 ( .a(stage_0[9][21]), .b(stage_0[9][22]), .cin(stage_0[9][23]), .cout(stage_1[10][7]), .s(stage_1[9][28]) );
FA FA_1_218 ( .a(stage_0[9][24]), .b(stage_0[9][25]), .cin(stage_0[9][26]), .cout(stage_1[10][8]), .s(stage_1[9][29]) );
FA FA_1_219 ( .a(stage_0[9][27]), .b(stage_0[9][28]), .cin(stage_0[9][29]), .cout(stage_1[10][9]), .s(stage_1[9][30]) );
FA FA_1_220 ( .a(stage_0[9][30]), .b(stage_0[9][31]), .cin(stage_0[9][32]), .cout(stage_1[10][10]), .s(stage_1[9][31]) );
FA FA_1_221 ( .a(stage_0[9][33]), .b(stage_0[9][34]), .cin(stage_0[9][35]), .cout(stage_1[10][11]), .s(stage_1[9][32]) );
FA FA_1_222 ( .a(stage_0[9][36]), .b(stage_0[9][37]), .cin(stage_0[9][38]), .cout(stage_1[10][12]), .s(stage_1[9][33]) );
FA FA_1_223 ( .a(stage_0[9][39]), .b(stage_0[9][40]), .cin(stage_0[9][41]), .cout(stage_1[10][13]), .s(stage_1[9][34]) );
FA FA_1_224 ( .a(stage_0[9][42]), .b(stage_0[9][43]), .cin(stage_0[9][44]), .cout(stage_1[10][14]), .s(stage_1[9][35]) );
FA FA_1_225 ( .a(stage_0[9][45]), .b(stage_0[9][46]), .cin(stage_0[9][47]), .cout(stage_1[10][15]), .s(stage_1[9][36]) );
FA FA_1_226 ( .a(stage_0[9][48]), .b(stage_0[9][49]), .cin(stage_0[9][50]), .cout(stage_1[10][16]), .s(stage_1[9][37]) );
FA FA_1_227 ( .a(stage_0[9][51]), .b(stage_0[9][52]), .cin(stage_0[9][53]), .cout(stage_1[10][17]), .s(stage_1[9][38]) );
FA FA_1_228 ( .a(stage_0[9][54]), .b(stage_0[9][55]), .cin(stage_0[9][56]), .cout(stage_1[10][18]), .s(stage_1[9][39]) );
FA FA_1_229 ( .a(stage_0[9][57]), .b(stage_0[9][58]), .cin(stage_0[9][59]), .cout(stage_1[10][19]), .s(stage_1[9][40]) );
FA FA_1_230 ( .a(stage_0[9][60]), .b(stage_0[9][61]), .cin(stage_0[9][62]), .cout(stage_1[10][20]), .s(stage_1[9][41]) );
assign stage_1[9][42] = stage_0[9][63];
FA FA_1_231 ( .a(stage_0[10][0]), .b(stage_0[10][1]), .cin(stage_0[10][2]), .cout(stage_1[11][0]), .s(stage_1[10][21]) );
FA FA_1_232 ( .a(stage_0[10][3]), .b(stage_0[10][4]), .cin(stage_0[10][5]), .cout(stage_1[11][1]), .s(stage_1[10][22]) );
FA FA_1_233 ( .a(stage_0[10][6]), .b(stage_0[10][7]), .cin(stage_0[10][8]), .cout(stage_1[11][2]), .s(stage_1[10][23]) );
FA FA_1_234 ( .a(stage_0[10][9]), .b(stage_0[10][10]), .cin(stage_0[10][11]), .cout(stage_1[11][3]), .s(stage_1[10][24]) );
FA FA_1_235 ( .a(stage_0[10][12]), .b(stage_0[10][13]), .cin(stage_0[10][14]), .cout(stage_1[11][4]), .s(stage_1[10][25]) );
FA FA_1_236 ( .a(stage_0[10][15]), .b(stage_0[10][16]), .cin(stage_0[10][17]), .cout(stage_1[11][5]), .s(stage_1[10][26]) );
FA FA_1_237 ( .a(stage_0[10][18]), .b(stage_0[10][19]), .cin(stage_0[10][20]), .cout(stage_1[11][6]), .s(stage_1[10][27]) );
FA FA_1_238 ( .a(stage_0[10][21]), .b(stage_0[10][22]), .cin(stage_0[10][23]), .cout(stage_1[11][7]), .s(stage_1[10][28]) );
FA FA_1_239 ( .a(stage_0[10][24]), .b(stage_0[10][25]), .cin(stage_0[10][26]), .cout(stage_1[11][8]), .s(stage_1[10][29]) );
FA FA_1_240 ( .a(stage_0[10][27]), .b(stage_0[10][28]), .cin(stage_0[10][29]), .cout(stage_1[11][9]), .s(stage_1[10][30]) );
FA FA_1_241 ( .a(stage_0[10][30]), .b(stage_0[10][31]), .cin(stage_0[10][32]), .cout(stage_1[11][10]), .s(stage_1[10][31]) );
FA FA_1_242 ( .a(stage_0[10][33]), .b(stage_0[10][34]), .cin(stage_0[10][35]), .cout(stage_1[11][11]), .s(stage_1[10][32]) );
FA FA_1_243 ( .a(stage_0[10][36]), .b(stage_0[10][37]), .cin(stage_0[10][38]), .cout(stage_1[11][12]), .s(stage_1[10][33]) );
FA FA_1_244 ( .a(stage_0[10][39]), .b(stage_0[10][40]), .cin(stage_0[10][41]), .cout(stage_1[11][13]), .s(stage_1[10][34]) );
FA FA_1_245 ( .a(stage_0[10][42]), .b(stage_0[10][43]), .cin(stage_0[10][44]), .cout(stage_1[11][14]), .s(stage_1[10][35]) );
FA FA_1_246 ( .a(stage_0[10][45]), .b(stage_0[10][46]), .cin(stage_0[10][47]), .cout(stage_1[11][15]), .s(stage_1[10][36]) );
FA FA_1_247 ( .a(stage_0[10][48]), .b(stage_0[10][49]), .cin(stage_0[10][50]), .cout(stage_1[11][16]), .s(stage_1[10][37]) );
FA FA_1_248 ( .a(stage_0[10][51]), .b(stage_0[10][52]), .cin(stage_0[10][53]), .cout(stage_1[11][17]), .s(stage_1[10][38]) );
FA FA_1_249 ( .a(stage_0[10][54]), .b(stage_0[10][55]), .cin(stage_0[10][56]), .cout(stage_1[11][18]), .s(stage_1[10][39]) );
FA FA_1_250 ( .a(stage_0[10][57]), .b(stage_0[10][58]), .cin(stage_0[10][59]), .cout(stage_1[11][19]), .s(stage_1[10][40]) );
FA FA_1_251 ( .a(stage_0[10][60]), .b(stage_0[10][61]), .cin(stage_0[10][62]), .cout(stage_1[11][20]), .s(stage_1[10][41]) );
assign stage_1[10][42] = stage_0[10][63];
FA FA_1_252 ( .a(stage_0[11][0]), .b(stage_0[11][1]), .cin(stage_0[11][2]), .cout(stage_1[12][0]), .s(stage_1[11][21]) );
FA FA_1_253 ( .a(stage_0[11][3]), .b(stage_0[11][4]), .cin(stage_0[11][5]), .cout(stage_1[12][1]), .s(stage_1[11][22]) );
FA FA_1_254 ( .a(stage_0[11][6]), .b(stage_0[11][7]), .cin(stage_0[11][8]), .cout(stage_1[12][2]), .s(stage_1[11][23]) );
FA FA_1_255 ( .a(stage_0[11][9]), .b(stage_0[11][10]), .cin(stage_0[11][11]), .cout(stage_1[12][3]), .s(stage_1[11][24]) );
FA FA_1_256 ( .a(stage_0[11][12]), .b(stage_0[11][13]), .cin(stage_0[11][14]), .cout(stage_1[12][4]), .s(stage_1[11][25]) );
FA FA_1_257 ( .a(stage_0[11][15]), .b(stage_0[11][16]), .cin(stage_0[11][17]), .cout(stage_1[12][5]), .s(stage_1[11][26]) );
FA FA_1_258 ( .a(stage_0[11][18]), .b(stage_0[11][19]), .cin(stage_0[11][20]), .cout(stage_1[12][6]), .s(stage_1[11][27]) );
FA FA_1_259 ( .a(stage_0[11][21]), .b(stage_0[11][22]), .cin(stage_0[11][23]), .cout(stage_1[12][7]), .s(stage_1[11][28]) );
FA FA_1_260 ( .a(stage_0[11][24]), .b(stage_0[11][25]), .cin(stage_0[11][26]), .cout(stage_1[12][8]), .s(stage_1[11][29]) );
FA FA_1_261 ( .a(stage_0[11][27]), .b(stage_0[11][28]), .cin(stage_0[11][29]), .cout(stage_1[12][9]), .s(stage_1[11][30]) );
FA FA_1_262 ( .a(stage_0[11][30]), .b(stage_0[11][31]), .cin(stage_0[11][32]), .cout(stage_1[12][10]), .s(stage_1[11][31]) );
FA FA_1_263 ( .a(stage_0[11][33]), .b(stage_0[11][34]), .cin(stage_0[11][35]), .cout(stage_1[12][11]), .s(stage_1[11][32]) );
FA FA_1_264 ( .a(stage_0[11][36]), .b(stage_0[11][37]), .cin(stage_0[11][38]), .cout(stage_1[12][12]), .s(stage_1[11][33]) );
FA FA_1_265 ( .a(stage_0[11][39]), .b(stage_0[11][40]), .cin(stage_0[11][41]), .cout(stage_1[12][13]), .s(stage_1[11][34]) );
FA FA_1_266 ( .a(stage_0[11][42]), .b(stage_0[11][43]), .cin(stage_0[11][44]), .cout(stage_1[12][14]), .s(stage_1[11][35]) );
FA FA_1_267 ( .a(stage_0[11][45]), .b(stage_0[11][46]), .cin(stage_0[11][47]), .cout(stage_1[12][15]), .s(stage_1[11][36]) );
FA FA_1_268 ( .a(stage_0[11][48]), .b(stage_0[11][49]), .cin(stage_0[11][50]), .cout(stage_1[12][16]), .s(stage_1[11][37]) );
FA FA_1_269 ( .a(stage_0[11][51]), .b(stage_0[11][52]), .cin(stage_0[11][53]), .cout(stage_1[12][17]), .s(stage_1[11][38]) );
FA FA_1_270 ( .a(stage_0[11][54]), .b(stage_0[11][55]), .cin(stage_0[11][56]), .cout(stage_1[12][18]), .s(stage_1[11][39]) );
FA FA_1_271 ( .a(stage_0[11][57]), .b(stage_0[11][58]), .cin(stage_0[11][59]), .cout(stage_1[12][19]), .s(stage_1[11][40]) );
FA FA_1_272 ( .a(stage_0[11][60]), .b(stage_0[11][61]), .cin(stage_0[11][62]), .cout(stage_1[12][20]), .s(stage_1[11][41]) );
assign stage_1[11][42] = stage_0[11][63];
FA FA_1_273 ( .a(stage_0[12][0]), .b(stage_0[12][1]), .cin(stage_0[12][2]), .cout(stage_1[13][0]), .s(stage_1[12][21]) );
FA FA_1_274 ( .a(stage_0[12][3]), .b(stage_0[12][4]), .cin(stage_0[12][5]), .cout(stage_1[13][1]), .s(stage_1[12][22]) );
FA FA_1_275 ( .a(stage_0[12][6]), .b(stage_0[12][7]), .cin(stage_0[12][8]), .cout(stage_1[13][2]), .s(stage_1[12][23]) );
FA FA_1_276 ( .a(stage_0[12][9]), .b(stage_0[12][10]), .cin(stage_0[12][11]), .cout(stage_1[13][3]), .s(stage_1[12][24]) );
FA FA_1_277 ( .a(stage_0[12][12]), .b(stage_0[12][13]), .cin(stage_0[12][14]), .cout(stage_1[13][4]), .s(stage_1[12][25]) );
FA FA_1_278 ( .a(stage_0[12][15]), .b(stage_0[12][16]), .cin(stage_0[12][17]), .cout(stage_1[13][5]), .s(stage_1[12][26]) );
FA FA_1_279 ( .a(stage_0[12][18]), .b(stage_0[12][19]), .cin(stage_0[12][20]), .cout(stage_1[13][6]), .s(stage_1[12][27]) );
FA FA_1_280 ( .a(stage_0[12][21]), .b(stage_0[12][22]), .cin(stage_0[12][23]), .cout(stage_1[13][7]), .s(stage_1[12][28]) );
FA FA_1_281 ( .a(stage_0[12][24]), .b(stage_0[12][25]), .cin(stage_0[12][26]), .cout(stage_1[13][8]), .s(stage_1[12][29]) );
FA FA_1_282 ( .a(stage_0[12][27]), .b(stage_0[12][28]), .cin(stage_0[12][29]), .cout(stage_1[13][9]), .s(stage_1[12][30]) );
FA FA_1_283 ( .a(stage_0[12][30]), .b(stage_0[12][31]), .cin(stage_0[12][32]), .cout(stage_1[13][10]), .s(stage_1[12][31]) );
FA FA_1_284 ( .a(stage_0[12][33]), .b(stage_0[12][34]), .cin(stage_0[12][35]), .cout(stage_1[13][11]), .s(stage_1[12][32]) );
FA FA_1_285 ( .a(stage_0[12][36]), .b(stage_0[12][37]), .cin(stage_0[12][38]), .cout(stage_1[13][12]), .s(stage_1[12][33]) );
FA FA_1_286 ( .a(stage_0[12][39]), .b(stage_0[12][40]), .cin(stage_0[12][41]), .cout(stage_1[13][13]), .s(stage_1[12][34]) );
FA FA_1_287 ( .a(stage_0[12][42]), .b(stage_0[12][43]), .cin(stage_0[12][44]), .cout(stage_1[13][14]), .s(stage_1[12][35]) );
FA FA_1_288 ( .a(stage_0[12][45]), .b(stage_0[12][46]), .cin(stage_0[12][47]), .cout(stage_1[13][15]), .s(stage_1[12][36]) );
FA FA_1_289 ( .a(stage_0[12][48]), .b(stage_0[12][49]), .cin(stage_0[12][50]), .cout(stage_1[13][16]), .s(stage_1[12][37]) );
FA FA_1_290 ( .a(stage_0[12][51]), .b(stage_0[12][52]), .cin(stage_0[12][53]), .cout(stage_1[13][17]), .s(stage_1[12][38]) );
FA FA_1_291 ( .a(stage_0[12][54]), .b(stage_0[12][55]), .cin(stage_0[12][56]), .cout(stage_1[13][18]), .s(stage_1[12][39]) );
FA FA_1_292 ( .a(stage_0[12][57]), .b(stage_0[12][58]), .cin(stage_0[12][59]), .cout(stage_1[13][19]), .s(stage_1[12][40]) );
FA FA_1_293 ( .a(stage_0[12][60]), .b(stage_0[12][61]), .cin(stage_0[12][62]), .cout(stage_1[13][20]), .s(stage_1[12][41]) );
assign stage_1[12][42] = stage_0[12][63];
FA FA_1_294 ( .a(stage_0[13][0]), .b(stage_0[13][1]), .cin(stage_0[13][2]), .cout(stage_1[14][0]), .s(stage_1[13][21]) );
FA FA_1_295 ( .a(stage_0[13][3]), .b(stage_0[13][4]), .cin(stage_0[13][5]), .cout(stage_1[14][1]), .s(stage_1[13][22]) );
FA FA_1_296 ( .a(stage_0[13][6]), .b(stage_0[13][7]), .cin(stage_0[13][8]), .cout(stage_1[14][2]), .s(stage_1[13][23]) );
FA FA_1_297 ( .a(stage_0[13][9]), .b(stage_0[13][10]), .cin(stage_0[13][11]), .cout(stage_1[14][3]), .s(stage_1[13][24]) );
FA FA_1_298 ( .a(stage_0[13][12]), .b(stage_0[13][13]), .cin(stage_0[13][14]), .cout(stage_1[14][4]), .s(stage_1[13][25]) );
FA FA_1_299 ( .a(stage_0[13][15]), .b(stage_0[13][16]), .cin(stage_0[13][17]), .cout(stage_1[14][5]), .s(stage_1[13][26]) );
FA FA_1_300 ( .a(stage_0[13][18]), .b(stage_0[13][19]), .cin(stage_0[13][20]), .cout(stage_1[14][6]), .s(stage_1[13][27]) );
FA FA_1_301 ( .a(stage_0[13][21]), .b(stage_0[13][22]), .cin(stage_0[13][23]), .cout(stage_1[14][7]), .s(stage_1[13][28]) );
FA FA_1_302 ( .a(stage_0[13][24]), .b(stage_0[13][25]), .cin(stage_0[13][26]), .cout(stage_1[14][8]), .s(stage_1[13][29]) );
FA FA_1_303 ( .a(stage_0[13][27]), .b(stage_0[13][28]), .cin(stage_0[13][29]), .cout(stage_1[14][9]), .s(stage_1[13][30]) );
FA FA_1_304 ( .a(stage_0[13][30]), .b(stage_0[13][31]), .cin(stage_0[13][32]), .cout(stage_1[14][10]), .s(stage_1[13][31]) );
FA FA_1_305 ( .a(stage_0[13][33]), .b(stage_0[13][34]), .cin(stage_0[13][35]), .cout(stage_1[14][11]), .s(stage_1[13][32]) );
FA FA_1_306 ( .a(stage_0[13][36]), .b(stage_0[13][37]), .cin(stage_0[13][38]), .cout(stage_1[14][12]), .s(stage_1[13][33]) );
FA FA_1_307 ( .a(stage_0[13][39]), .b(stage_0[13][40]), .cin(stage_0[13][41]), .cout(stage_1[14][13]), .s(stage_1[13][34]) );
FA FA_1_308 ( .a(stage_0[13][42]), .b(stage_0[13][43]), .cin(stage_0[13][44]), .cout(stage_1[14][14]), .s(stage_1[13][35]) );
FA FA_1_309 ( .a(stage_0[13][45]), .b(stage_0[13][46]), .cin(stage_0[13][47]), .cout(stage_1[14][15]), .s(stage_1[13][36]) );
FA FA_1_310 ( .a(stage_0[13][48]), .b(stage_0[13][49]), .cin(stage_0[13][50]), .cout(stage_1[14][16]), .s(stage_1[13][37]) );
FA FA_1_311 ( .a(stage_0[13][51]), .b(stage_0[13][52]), .cin(stage_0[13][53]), .cout(stage_1[14][17]), .s(stage_1[13][38]) );
FA FA_1_312 ( .a(stage_0[13][54]), .b(stage_0[13][55]), .cin(stage_0[13][56]), .cout(stage_1[14][18]), .s(stage_1[13][39]) );
FA FA_1_313 ( .a(stage_0[13][57]), .b(stage_0[13][58]), .cin(stage_0[13][59]), .cout(stage_1[14][19]), .s(stage_1[13][40]) );
FA FA_1_314 ( .a(stage_0[13][60]), .b(stage_0[13][61]), .cin(stage_0[13][62]), .cout(stage_1[14][20]), .s(stage_1[13][41]) );
assign stage_1[13][42] = stage_0[13][63];
FA FA_1_315 ( .a(stage_0[14][0]), .b(stage_0[14][1]), .cin(stage_0[14][2]), .cout(stage_1[15][0]), .s(stage_1[14][21]) );
FA FA_1_316 ( .a(stage_0[14][3]), .b(stage_0[14][4]), .cin(stage_0[14][5]), .cout(stage_1[15][1]), .s(stage_1[14][22]) );
FA FA_1_317 ( .a(stage_0[14][6]), .b(stage_0[14][7]), .cin(stage_0[14][8]), .cout(stage_1[15][2]), .s(stage_1[14][23]) );
FA FA_1_318 ( .a(stage_0[14][9]), .b(stage_0[14][10]), .cin(stage_0[14][11]), .cout(stage_1[15][3]), .s(stage_1[14][24]) );
FA FA_1_319 ( .a(stage_0[14][12]), .b(stage_0[14][13]), .cin(stage_0[14][14]), .cout(stage_1[15][4]), .s(stage_1[14][25]) );
FA FA_1_320 ( .a(stage_0[14][15]), .b(stage_0[14][16]), .cin(stage_0[14][17]), .cout(stage_1[15][5]), .s(stage_1[14][26]) );
FA FA_1_321 ( .a(stage_0[14][18]), .b(stage_0[14][19]), .cin(stage_0[14][20]), .cout(stage_1[15][6]), .s(stage_1[14][27]) );
FA FA_1_322 ( .a(stage_0[14][21]), .b(stage_0[14][22]), .cin(stage_0[14][23]), .cout(stage_1[15][7]), .s(stage_1[14][28]) );
FA FA_1_323 ( .a(stage_0[14][24]), .b(stage_0[14][25]), .cin(stage_0[14][26]), .cout(stage_1[15][8]), .s(stage_1[14][29]) );
FA FA_1_324 ( .a(stage_0[14][27]), .b(stage_0[14][28]), .cin(stage_0[14][29]), .cout(stage_1[15][9]), .s(stage_1[14][30]) );
FA FA_1_325 ( .a(stage_0[14][30]), .b(stage_0[14][31]), .cin(stage_0[14][32]), .cout(stage_1[15][10]), .s(stage_1[14][31]) );
FA FA_1_326 ( .a(stage_0[14][33]), .b(stage_0[14][34]), .cin(stage_0[14][35]), .cout(stage_1[15][11]), .s(stage_1[14][32]) );
FA FA_1_327 ( .a(stage_0[14][36]), .b(stage_0[14][37]), .cin(stage_0[14][38]), .cout(stage_1[15][12]), .s(stage_1[14][33]) );
FA FA_1_328 ( .a(stage_0[14][39]), .b(stage_0[14][40]), .cin(stage_0[14][41]), .cout(stage_1[15][13]), .s(stage_1[14][34]) );
FA FA_1_329 ( .a(stage_0[14][42]), .b(stage_0[14][43]), .cin(stage_0[14][44]), .cout(stage_1[15][14]), .s(stage_1[14][35]) );
FA FA_1_330 ( .a(stage_0[14][45]), .b(stage_0[14][46]), .cin(stage_0[14][47]), .cout(stage_1[15][15]), .s(stage_1[14][36]) );
FA FA_1_331 ( .a(stage_0[14][48]), .b(stage_0[14][49]), .cin(stage_0[14][50]), .cout(stage_1[15][16]), .s(stage_1[14][37]) );
FA FA_1_332 ( .a(stage_0[14][51]), .b(stage_0[14][52]), .cin(stage_0[14][53]), .cout(stage_1[15][17]), .s(stage_1[14][38]) );
FA FA_1_333 ( .a(stage_0[14][54]), .b(stage_0[14][55]), .cin(stage_0[14][56]), .cout(stage_1[15][18]), .s(stage_1[14][39]) );
FA FA_1_334 ( .a(stage_0[14][57]), .b(stage_0[14][58]), .cin(stage_0[14][59]), .cout(stage_1[15][19]), .s(stage_1[14][40]) );
FA FA_1_335 ( .a(stage_0[14][60]), .b(stage_0[14][61]), .cin(stage_0[14][62]), .cout(stage_1[15][20]), .s(stage_1[14][41]) );
assign stage_1[14][42] = stage_0[14][63];
FA FA_1_336 ( .a(stage_0[15][0]), .b(stage_0[15][1]), .cin(stage_0[15][2]), .cout(stage_1[16][0]), .s(stage_1[15][21]) );
FA FA_1_337 ( .a(stage_0[15][3]), .b(stage_0[15][4]), .cin(stage_0[15][5]), .cout(stage_1[16][1]), .s(stage_1[15][22]) );
FA FA_1_338 ( .a(stage_0[15][6]), .b(stage_0[15][7]), .cin(stage_0[15][8]), .cout(stage_1[16][2]), .s(stage_1[15][23]) );
FA FA_1_339 ( .a(stage_0[15][9]), .b(stage_0[15][10]), .cin(stage_0[15][11]), .cout(stage_1[16][3]), .s(stage_1[15][24]) );
FA FA_1_340 ( .a(stage_0[15][12]), .b(stage_0[15][13]), .cin(stage_0[15][14]), .cout(stage_1[16][4]), .s(stage_1[15][25]) );
FA FA_1_341 ( .a(stage_0[15][15]), .b(stage_0[15][16]), .cin(stage_0[15][17]), .cout(stage_1[16][5]), .s(stage_1[15][26]) );
FA FA_1_342 ( .a(stage_0[15][18]), .b(stage_0[15][19]), .cin(stage_0[15][20]), .cout(stage_1[16][6]), .s(stage_1[15][27]) );
FA FA_1_343 ( .a(stage_0[15][21]), .b(stage_0[15][22]), .cin(stage_0[15][23]), .cout(stage_1[16][7]), .s(stage_1[15][28]) );
FA FA_1_344 ( .a(stage_0[15][24]), .b(stage_0[15][25]), .cin(stage_0[15][26]), .cout(stage_1[16][8]), .s(stage_1[15][29]) );
FA FA_1_345 ( .a(stage_0[15][27]), .b(stage_0[15][28]), .cin(stage_0[15][29]), .cout(stage_1[16][9]), .s(stage_1[15][30]) );
FA FA_1_346 ( .a(stage_0[15][30]), .b(stage_0[15][31]), .cin(stage_0[15][32]), .cout(stage_1[16][10]), .s(stage_1[15][31]) );
FA FA_1_347 ( .a(stage_0[15][33]), .b(stage_0[15][34]), .cin(stage_0[15][35]), .cout(stage_1[16][11]), .s(stage_1[15][32]) );
FA FA_1_348 ( .a(stage_0[15][36]), .b(stage_0[15][37]), .cin(stage_0[15][38]), .cout(stage_1[16][12]), .s(stage_1[15][33]) );
FA FA_1_349 ( .a(stage_0[15][39]), .b(stage_0[15][40]), .cin(stage_0[15][41]), .cout(stage_1[16][13]), .s(stage_1[15][34]) );
FA FA_1_350 ( .a(stage_0[15][42]), .b(stage_0[15][43]), .cin(stage_0[15][44]), .cout(stage_1[16][14]), .s(stage_1[15][35]) );
FA FA_1_351 ( .a(stage_0[15][45]), .b(stage_0[15][46]), .cin(stage_0[15][47]), .cout(stage_1[16][15]), .s(stage_1[15][36]) );
FA FA_1_352 ( .a(stage_0[15][48]), .b(stage_0[15][49]), .cin(stage_0[15][50]), .cout(stage_1[16][16]), .s(stage_1[15][37]) );
FA FA_1_353 ( .a(stage_0[15][51]), .b(stage_0[15][52]), .cin(stage_0[15][53]), .cout(stage_1[16][17]), .s(stage_1[15][38]) );
FA FA_1_354 ( .a(stage_0[15][54]), .b(stage_0[15][55]), .cin(stage_0[15][56]), .cout(stage_1[16][18]), .s(stage_1[15][39]) );
FA FA_1_355 ( .a(stage_0[15][57]), .b(stage_0[15][58]), .cin(stage_0[15][59]), .cout(stage_1[16][19]), .s(stage_1[15][40]) );
FA FA_1_356 ( .a(stage_0[15][60]), .b(stage_0[15][61]), .cin(stage_0[15][62]), .cout(stage_1[16][20]), .s(stage_1[15][41]) );
assign stage_1[15][42] = stage_0[15][63];

wire stage_2 [`NBIT+2:0][`NDATA*2:0];
FA FA_2_0 ( .a(stage_1[0][0]), .b(stage_1[0][1]), .cin(stage_1[0][2]), .cout(stage_2[1][0]), .s(stage_2[0][0]) );
FA FA_2_1 ( .a(stage_1[0][3]), .b(stage_1[0][4]), .cin(stage_1[0][5]), .cout(stage_2[1][1]), .s(stage_2[0][1]) );
FA FA_2_2 ( .a(stage_1[0][6]), .b(stage_1[0][7]), .cin(stage_1[0][8]), .cout(stage_2[1][2]), .s(stage_2[0][2]) );
FA FA_2_3 ( .a(stage_1[0][9]), .b(stage_1[0][10]), .cin(stage_1[0][11]), .cout(stage_2[1][3]), .s(stage_2[0][3]) );
FA FA_2_4 ( .a(stage_1[0][12]), .b(stage_1[0][13]), .cin(stage_1[0][14]), .cout(stage_2[1][4]), .s(stage_2[0][4]) );
FA FA_2_5 ( .a(stage_1[0][15]), .b(stage_1[0][16]), .cin(stage_1[0][17]), .cout(stage_2[1][5]), .s(stage_2[0][5]) );
FA FA_2_6 ( .a(stage_1[0][18]), .b(stage_1[0][19]), .cin(stage_1[0][20]), .cout(stage_2[1][6]), .s(stage_2[0][6]) );
FA FA_2_7 ( .a(stage_1[0][21]), .b(stage_1[0][22]), .cin(stage_1[0][23]), .cout(stage_2[1][7]), .s(stage_2[0][7]) );
FA FA_2_8 ( .a(stage_1[0][24]), .b(stage_1[0][25]), .cin(stage_1[0][26]), .cout(stage_2[1][8]), .s(stage_2[0][8]) );
FA FA_2_9 ( .a(stage_1[0][27]), .b(stage_1[0][28]), .cin(stage_1[0][29]), .cout(stage_2[1][9]), .s(stage_2[0][9]) );
FA FA_2_10 ( .a(stage_1[0][30]), .b(stage_1[0][31]), .cin(stage_1[0][32]), .cout(stage_2[1][10]), .s(stage_2[0][10]) );
FA FA_2_11 ( .a(stage_1[0][33]), .b(stage_1[0][34]), .cin(stage_1[0][35]), .cout(stage_2[1][11]), .s(stage_2[0][11]) );
FA FA_2_12 ( .a(stage_1[0][36]), .b(stage_1[0][37]), .cin(stage_1[0][38]), .cout(stage_2[1][12]), .s(stage_2[0][12]) );
FA FA_2_13 ( .a(stage_1[0][39]), .b(stage_1[0][40]), .cin(stage_1[0][41]), .cout(stage_2[1][13]), .s(stage_2[0][13]) );
assign stage_2[0][14] = stage_1[0][42];
FA FA_2_14 ( .a(stage_1[1][0]), .b(stage_1[1][1]), .cin(stage_1[1][2]), .cout(stage_2[2][0]), .s(stage_2[1][14]) );
FA FA_2_15 ( .a(stage_1[1][3]), .b(stage_1[1][4]), .cin(stage_1[1][5]), .cout(stage_2[2][1]), .s(stage_2[1][15]) );
FA FA_2_16 ( .a(stage_1[1][6]), .b(stage_1[1][7]), .cin(stage_1[1][8]), .cout(stage_2[2][2]), .s(stage_2[1][16]) );
FA FA_2_17 ( .a(stage_1[1][9]), .b(stage_1[1][10]), .cin(stage_1[1][11]), .cout(stage_2[2][3]), .s(stage_2[1][17]) );
FA FA_2_18 ( .a(stage_1[1][12]), .b(stage_1[1][13]), .cin(stage_1[1][14]), .cout(stage_2[2][4]), .s(stage_2[1][18]) );
FA FA_2_19 ( .a(stage_1[1][15]), .b(stage_1[1][16]), .cin(stage_1[1][17]), .cout(stage_2[2][5]), .s(stage_2[1][19]) );
FA FA_2_20 ( .a(stage_1[1][18]), .b(stage_1[1][19]), .cin(stage_1[1][20]), .cout(stage_2[2][6]), .s(stage_2[1][20]) );
FA FA_2_21 ( .a(stage_1[1][21]), .b(stage_1[1][22]), .cin(stage_1[1][23]), .cout(stage_2[2][7]), .s(stage_2[1][21]) );
FA FA_2_22 ( .a(stage_1[1][24]), .b(stage_1[1][25]), .cin(stage_1[1][26]), .cout(stage_2[2][8]), .s(stage_2[1][22]) );
FA FA_2_23 ( .a(stage_1[1][27]), .b(stage_1[1][28]), .cin(stage_1[1][29]), .cout(stage_2[2][9]), .s(stage_2[1][23]) );
FA FA_2_24 ( .a(stage_1[1][30]), .b(stage_1[1][31]), .cin(stage_1[1][32]), .cout(stage_2[2][10]), .s(stage_2[1][24]) );
FA FA_2_25 ( .a(stage_1[1][33]), .b(stage_1[1][34]), .cin(stage_1[1][35]), .cout(stage_2[2][11]), .s(stage_2[1][25]) );
FA FA_2_26 ( .a(stage_1[1][36]), .b(stage_1[1][37]), .cin(stage_1[1][38]), .cout(stage_2[2][12]), .s(stage_2[1][26]) );
FA FA_2_27 ( .a(stage_1[1][39]), .b(stage_1[1][40]), .cin(stage_1[1][41]), .cout(stage_2[2][13]), .s(stage_2[1][27]) );
FA FA_2_28 ( .a(stage_1[1][42]), .b(stage_1[1][43]), .cin(stage_1[1][44]), .cout(stage_2[2][14]), .s(stage_2[1][28]) );
FA FA_2_29 ( .a(stage_1[1][45]), .b(stage_1[1][46]), .cin(stage_1[1][47]), .cout(stage_2[2][15]), .s(stage_2[1][29]) );
FA FA_2_30 ( .a(stage_1[1][48]), .b(stage_1[1][49]), .cin(stage_1[1][50]), .cout(stage_2[2][16]), .s(stage_2[1][30]) );
FA FA_2_31 ( .a(stage_1[1][51]), .b(stage_1[1][52]), .cin(stage_1[1][53]), .cout(stage_2[2][17]), .s(stage_2[1][31]) );
FA FA_2_32 ( .a(stage_1[1][54]), .b(stage_1[1][55]), .cin(stage_1[1][56]), .cout(stage_2[2][18]), .s(stage_2[1][32]) );
FA FA_2_33 ( .a(stage_1[1][57]), .b(stage_1[1][58]), .cin(stage_1[1][59]), .cout(stage_2[2][19]), .s(stage_2[1][33]) );
FA FA_2_34 ( .a(stage_1[1][60]), .b(stage_1[1][61]), .cin(stage_1[1][62]), .cout(stage_2[2][20]), .s(stage_2[1][34]) );
HA HA_2_0 ( .a(stage_1[1][63]), .b(stage_1[1][64]), .cout(stage_2[2][21]), .s(stage_2[1][35]) );
FA FA_2_35 ( .a(stage_1[2][0]), .b(stage_1[2][1]), .cin(stage_1[2][2]), .cout(stage_2[3][0]), .s(stage_2[2][22]) );
FA FA_2_36 ( .a(stage_1[2][3]), .b(stage_1[2][4]), .cin(stage_1[2][5]), .cout(stage_2[3][1]), .s(stage_2[2][23]) );
FA FA_2_37 ( .a(stage_1[2][6]), .b(stage_1[2][7]), .cin(stage_1[2][8]), .cout(stage_2[3][2]), .s(stage_2[2][24]) );
FA FA_2_38 ( .a(stage_1[2][9]), .b(stage_1[2][10]), .cin(stage_1[2][11]), .cout(stage_2[3][3]), .s(stage_2[2][25]) );
FA FA_2_39 ( .a(stage_1[2][12]), .b(stage_1[2][13]), .cin(stage_1[2][14]), .cout(stage_2[3][4]), .s(stage_2[2][26]) );
FA FA_2_40 ( .a(stage_1[2][15]), .b(stage_1[2][16]), .cin(stage_1[2][17]), .cout(stage_2[3][5]), .s(stage_2[2][27]) );
FA FA_2_41 ( .a(stage_1[2][18]), .b(stage_1[2][19]), .cin(stage_1[2][20]), .cout(stage_2[3][6]), .s(stage_2[2][28]) );
FA FA_2_42 ( .a(stage_1[2][21]), .b(stage_1[2][22]), .cin(stage_1[2][23]), .cout(stage_2[3][7]), .s(stage_2[2][29]) );
FA FA_2_43 ( .a(stage_1[2][24]), .b(stage_1[2][25]), .cin(stage_1[2][26]), .cout(stage_2[3][8]), .s(stage_2[2][30]) );
FA FA_2_44 ( .a(stage_1[2][27]), .b(stage_1[2][28]), .cin(stage_1[2][29]), .cout(stage_2[3][9]), .s(stage_2[2][31]) );
FA FA_2_45 ( .a(stage_1[2][30]), .b(stage_1[2][31]), .cin(stage_1[2][32]), .cout(stage_2[3][10]), .s(stage_2[2][32]) );
FA FA_2_46 ( .a(stage_1[2][33]), .b(stage_1[2][34]), .cin(stage_1[2][35]), .cout(stage_2[3][11]), .s(stage_2[2][33]) );
FA FA_2_47 ( .a(stage_1[2][36]), .b(stage_1[2][37]), .cin(stage_1[2][38]), .cout(stage_2[3][12]), .s(stage_2[2][34]) );
FA FA_2_48 ( .a(stage_1[2][39]), .b(stage_1[2][40]), .cin(stage_1[2][41]), .cout(stage_2[3][13]), .s(stage_2[2][35]) );
assign stage_2[2][36] = stage_1[2][42];
FA FA_2_49 ( .a(stage_1[3][0]), .b(stage_1[3][1]), .cin(stage_1[3][2]), .cout(stage_2[4][0]), .s(stage_2[3][14]) );
FA FA_2_50 ( .a(stage_1[3][3]), .b(stage_1[3][4]), .cin(stage_1[3][5]), .cout(stage_2[4][1]), .s(stage_2[3][15]) );
FA FA_2_51 ( .a(stage_1[3][6]), .b(stage_1[3][7]), .cin(stage_1[3][8]), .cout(stage_2[4][2]), .s(stage_2[3][16]) );
FA FA_2_52 ( .a(stage_1[3][9]), .b(stage_1[3][10]), .cin(stage_1[3][11]), .cout(stage_2[4][3]), .s(stage_2[3][17]) );
FA FA_2_53 ( .a(stage_1[3][12]), .b(stage_1[3][13]), .cin(stage_1[3][14]), .cout(stage_2[4][4]), .s(stage_2[3][18]) );
FA FA_2_54 ( .a(stage_1[3][15]), .b(stage_1[3][16]), .cin(stage_1[3][17]), .cout(stage_2[4][5]), .s(stage_2[3][19]) );
FA FA_2_55 ( .a(stage_1[3][18]), .b(stage_1[3][19]), .cin(stage_1[3][20]), .cout(stage_2[4][6]), .s(stage_2[3][20]) );
FA FA_2_56 ( .a(stage_1[3][21]), .b(stage_1[3][22]), .cin(stage_1[3][23]), .cout(stage_2[4][7]), .s(stage_2[3][21]) );
FA FA_2_57 ( .a(stage_1[3][24]), .b(stage_1[3][25]), .cin(stage_1[3][26]), .cout(stage_2[4][8]), .s(stage_2[3][22]) );
FA FA_2_58 ( .a(stage_1[3][27]), .b(stage_1[3][28]), .cin(stage_1[3][29]), .cout(stage_2[4][9]), .s(stage_2[3][23]) );
FA FA_2_59 ( .a(stage_1[3][30]), .b(stage_1[3][31]), .cin(stage_1[3][32]), .cout(stage_2[4][10]), .s(stage_2[3][24]) );
FA FA_2_60 ( .a(stage_1[3][33]), .b(stage_1[3][34]), .cin(stage_1[3][35]), .cout(stage_2[4][11]), .s(stage_2[3][25]) );
FA FA_2_61 ( .a(stage_1[3][36]), .b(stage_1[3][37]), .cin(stage_1[3][38]), .cout(stage_2[4][12]), .s(stage_2[3][26]) );
FA FA_2_62 ( .a(stage_1[3][39]), .b(stage_1[3][40]), .cin(stage_1[3][41]), .cout(stage_2[4][13]), .s(stage_2[3][27]) );
assign stage_2[3][28] = stage_1[3][42];
FA FA_2_63 ( .a(stage_1[4][0]), .b(stage_1[4][1]), .cin(stage_1[4][2]), .cout(stage_2[5][0]), .s(stage_2[4][14]) );
FA FA_2_64 ( .a(stage_1[4][3]), .b(stage_1[4][4]), .cin(stage_1[4][5]), .cout(stage_2[5][1]), .s(stage_2[4][15]) );
FA FA_2_65 ( .a(stage_1[4][6]), .b(stage_1[4][7]), .cin(stage_1[4][8]), .cout(stage_2[5][2]), .s(stage_2[4][16]) );
FA FA_2_66 ( .a(stage_1[4][9]), .b(stage_1[4][10]), .cin(stage_1[4][11]), .cout(stage_2[5][3]), .s(stage_2[4][17]) );
FA FA_2_67 ( .a(stage_1[4][12]), .b(stage_1[4][13]), .cin(stage_1[4][14]), .cout(stage_2[5][4]), .s(stage_2[4][18]) );
FA FA_2_68 ( .a(stage_1[4][15]), .b(stage_1[4][16]), .cin(stage_1[4][17]), .cout(stage_2[5][5]), .s(stage_2[4][19]) );
FA FA_2_69 ( .a(stage_1[4][18]), .b(stage_1[4][19]), .cin(stage_1[4][20]), .cout(stage_2[5][6]), .s(stage_2[4][20]) );
FA FA_2_70 ( .a(stage_1[4][21]), .b(stage_1[4][22]), .cin(stage_1[4][23]), .cout(stage_2[5][7]), .s(stage_2[4][21]) );
FA FA_2_71 ( .a(stage_1[4][24]), .b(stage_1[4][25]), .cin(stage_1[4][26]), .cout(stage_2[5][8]), .s(stage_2[4][22]) );
FA FA_2_72 ( .a(stage_1[4][27]), .b(stage_1[4][28]), .cin(stage_1[4][29]), .cout(stage_2[5][9]), .s(stage_2[4][23]) );
FA FA_2_73 ( .a(stage_1[4][30]), .b(stage_1[4][31]), .cin(stage_1[4][32]), .cout(stage_2[5][10]), .s(stage_2[4][24]) );
FA FA_2_74 ( .a(stage_1[4][33]), .b(stage_1[4][34]), .cin(stage_1[4][35]), .cout(stage_2[5][11]), .s(stage_2[4][25]) );
FA FA_2_75 ( .a(stage_1[4][36]), .b(stage_1[4][37]), .cin(stage_1[4][38]), .cout(stage_2[5][12]), .s(stage_2[4][26]) );
FA FA_2_76 ( .a(stage_1[4][39]), .b(stage_1[4][40]), .cin(stage_1[4][41]), .cout(stage_2[5][13]), .s(stage_2[4][27]) );
assign stage_2[4][28] = stage_1[4][42];
FA FA_2_77 ( .a(stage_1[5][0]), .b(stage_1[5][1]), .cin(stage_1[5][2]), .cout(stage_2[6][0]), .s(stage_2[5][14]) );
FA FA_2_78 ( .a(stage_1[5][3]), .b(stage_1[5][4]), .cin(stage_1[5][5]), .cout(stage_2[6][1]), .s(stage_2[5][15]) );
FA FA_2_79 ( .a(stage_1[5][6]), .b(stage_1[5][7]), .cin(stage_1[5][8]), .cout(stage_2[6][2]), .s(stage_2[5][16]) );
FA FA_2_80 ( .a(stage_1[5][9]), .b(stage_1[5][10]), .cin(stage_1[5][11]), .cout(stage_2[6][3]), .s(stage_2[5][17]) );
FA FA_2_81 ( .a(stage_1[5][12]), .b(stage_1[5][13]), .cin(stage_1[5][14]), .cout(stage_2[6][4]), .s(stage_2[5][18]) );
FA FA_2_82 ( .a(stage_1[5][15]), .b(stage_1[5][16]), .cin(stage_1[5][17]), .cout(stage_2[6][5]), .s(stage_2[5][19]) );
FA FA_2_83 ( .a(stage_1[5][18]), .b(stage_1[5][19]), .cin(stage_1[5][20]), .cout(stage_2[6][6]), .s(stage_2[5][20]) );
FA FA_2_84 ( .a(stage_1[5][21]), .b(stage_1[5][22]), .cin(stage_1[5][23]), .cout(stage_2[6][7]), .s(stage_2[5][21]) );
FA FA_2_85 ( .a(stage_1[5][24]), .b(stage_1[5][25]), .cin(stage_1[5][26]), .cout(stage_2[6][8]), .s(stage_2[5][22]) );
FA FA_2_86 ( .a(stage_1[5][27]), .b(stage_1[5][28]), .cin(stage_1[5][29]), .cout(stage_2[6][9]), .s(stage_2[5][23]) );
FA FA_2_87 ( .a(stage_1[5][30]), .b(stage_1[5][31]), .cin(stage_1[5][32]), .cout(stage_2[6][10]), .s(stage_2[5][24]) );
FA FA_2_88 ( .a(stage_1[5][33]), .b(stage_1[5][34]), .cin(stage_1[5][35]), .cout(stage_2[6][11]), .s(stage_2[5][25]) );
FA FA_2_89 ( .a(stage_1[5][36]), .b(stage_1[5][37]), .cin(stage_1[5][38]), .cout(stage_2[6][12]), .s(stage_2[5][26]) );
FA FA_2_90 ( .a(stage_1[5][39]), .b(stage_1[5][40]), .cin(stage_1[5][41]), .cout(stage_2[6][13]), .s(stage_2[5][27]) );
assign stage_2[5][28] = stage_1[5][42];
FA FA_2_91 ( .a(stage_1[6][0]), .b(stage_1[6][1]), .cin(stage_1[6][2]), .cout(stage_2[7][0]), .s(stage_2[6][14]) );
FA FA_2_92 ( .a(stage_1[6][3]), .b(stage_1[6][4]), .cin(stage_1[6][5]), .cout(stage_2[7][1]), .s(stage_2[6][15]) );
FA FA_2_93 ( .a(stage_1[6][6]), .b(stage_1[6][7]), .cin(stage_1[6][8]), .cout(stage_2[7][2]), .s(stage_2[6][16]) );
FA FA_2_94 ( .a(stage_1[6][9]), .b(stage_1[6][10]), .cin(stage_1[6][11]), .cout(stage_2[7][3]), .s(stage_2[6][17]) );
FA FA_2_95 ( .a(stage_1[6][12]), .b(stage_1[6][13]), .cin(stage_1[6][14]), .cout(stage_2[7][4]), .s(stage_2[6][18]) );
FA FA_2_96 ( .a(stage_1[6][15]), .b(stage_1[6][16]), .cin(stage_1[6][17]), .cout(stage_2[7][5]), .s(stage_2[6][19]) );
FA FA_2_97 ( .a(stage_1[6][18]), .b(stage_1[6][19]), .cin(stage_1[6][20]), .cout(stage_2[7][6]), .s(stage_2[6][20]) );
FA FA_2_98 ( .a(stage_1[6][21]), .b(stage_1[6][22]), .cin(stage_1[6][23]), .cout(stage_2[7][7]), .s(stage_2[6][21]) );
FA FA_2_99 ( .a(stage_1[6][24]), .b(stage_1[6][25]), .cin(stage_1[6][26]), .cout(stage_2[7][8]), .s(stage_2[6][22]) );
FA FA_2_100 ( .a(stage_1[6][27]), .b(stage_1[6][28]), .cin(stage_1[6][29]), .cout(stage_2[7][9]), .s(stage_2[6][23]) );
FA FA_2_101 ( .a(stage_1[6][30]), .b(stage_1[6][31]), .cin(stage_1[6][32]), .cout(stage_2[7][10]), .s(stage_2[6][24]) );
FA FA_2_102 ( .a(stage_1[6][33]), .b(stage_1[6][34]), .cin(stage_1[6][35]), .cout(stage_2[7][11]), .s(stage_2[6][25]) );
FA FA_2_103 ( .a(stage_1[6][36]), .b(stage_1[6][37]), .cin(stage_1[6][38]), .cout(stage_2[7][12]), .s(stage_2[6][26]) );
FA FA_2_104 ( .a(stage_1[6][39]), .b(stage_1[6][40]), .cin(stage_1[6][41]), .cout(stage_2[7][13]), .s(stage_2[6][27]) );
assign stage_2[6][28] = stage_1[6][42];
FA FA_2_105 ( .a(stage_1[7][0]), .b(stage_1[7][1]), .cin(stage_1[7][2]), .cout(stage_2[8][0]), .s(stage_2[7][14]) );
FA FA_2_106 ( .a(stage_1[7][3]), .b(stage_1[7][4]), .cin(stage_1[7][5]), .cout(stage_2[8][1]), .s(stage_2[7][15]) );
FA FA_2_107 ( .a(stage_1[7][6]), .b(stage_1[7][7]), .cin(stage_1[7][8]), .cout(stage_2[8][2]), .s(stage_2[7][16]) );
FA FA_2_108 ( .a(stage_1[7][9]), .b(stage_1[7][10]), .cin(stage_1[7][11]), .cout(stage_2[8][3]), .s(stage_2[7][17]) );
FA FA_2_109 ( .a(stage_1[7][12]), .b(stage_1[7][13]), .cin(stage_1[7][14]), .cout(stage_2[8][4]), .s(stage_2[7][18]) );
FA FA_2_110 ( .a(stage_1[7][15]), .b(stage_1[7][16]), .cin(stage_1[7][17]), .cout(stage_2[8][5]), .s(stage_2[7][19]) );
FA FA_2_111 ( .a(stage_1[7][18]), .b(stage_1[7][19]), .cin(stage_1[7][20]), .cout(stage_2[8][6]), .s(stage_2[7][20]) );
FA FA_2_112 ( .a(stage_1[7][21]), .b(stage_1[7][22]), .cin(stage_1[7][23]), .cout(stage_2[8][7]), .s(stage_2[7][21]) );
FA FA_2_113 ( .a(stage_1[7][24]), .b(stage_1[7][25]), .cin(stage_1[7][26]), .cout(stage_2[8][8]), .s(stage_2[7][22]) );
FA FA_2_114 ( .a(stage_1[7][27]), .b(stage_1[7][28]), .cin(stage_1[7][29]), .cout(stage_2[8][9]), .s(stage_2[7][23]) );
FA FA_2_115 ( .a(stage_1[7][30]), .b(stage_1[7][31]), .cin(stage_1[7][32]), .cout(stage_2[8][10]), .s(stage_2[7][24]) );
FA FA_2_116 ( .a(stage_1[7][33]), .b(stage_1[7][34]), .cin(stage_1[7][35]), .cout(stage_2[8][11]), .s(stage_2[7][25]) );
FA FA_2_117 ( .a(stage_1[7][36]), .b(stage_1[7][37]), .cin(stage_1[7][38]), .cout(stage_2[8][12]), .s(stage_2[7][26]) );
FA FA_2_118 ( .a(stage_1[7][39]), .b(stage_1[7][40]), .cin(stage_1[7][41]), .cout(stage_2[8][13]), .s(stage_2[7][27]) );
assign stage_2[7][28] = stage_1[7][42];
FA FA_2_119 ( .a(stage_1[8][0]), .b(stage_1[8][1]), .cin(stage_1[8][2]), .cout(stage_2[9][0]), .s(stage_2[8][14]) );
FA FA_2_120 ( .a(stage_1[8][3]), .b(stage_1[8][4]), .cin(stage_1[8][5]), .cout(stage_2[9][1]), .s(stage_2[8][15]) );
FA FA_2_121 ( .a(stage_1[8][6]), .b(stage_1[8][7]), .cin(stage_1[8][8]), .cout(stage_2[9][2]), .s(stage_2[8][16]) );
FA FA_2_122 ( .a(stage_1[8][9]), .b(stage_1[8][10]), .cin(stage_1[8][11]), .cout(stage_2[9][3]), .s(stage_2[8][17]) );
FA FA_2_123 ( .a(stage_1[8][12]), .b(stage_1[8][13]), .cin(stage_1[8][14]), .cout(stage_2[9][4]), .s(stage_2[8][18]) );
FA FA_2_124 ( .a(stage_1[8][15]), .b(stage_1[8][16]), .cin(stage_1[8][17]), .cout(stage_2[9][5]), .s(stage_2[8][19]) );
FA FA_2_125 ( .a(stage_1[8][18]), .b(stage_1[8][19]), .cin(stage_1[8][20]), .cout(stage_2[9][6]), .s(stage_2[8][20]) );
FA FA_2_126 ( .a(stage_1[8][21]), .b(stage_1[8][22]), .cin(stage_1[8][23]), .cout(stage_2[9][7]), .s(stage_2[8][21]) );
FA FA_2_127 ( .a(stage_1[8][24]), .b(stage_1[8][25]), .cin(stage_1[8][26]), .cout(stage_2[9][8]), .s(stage_2[8][22]) );
FA FA_2_128 ( .a(stage_1[8][27]), .b(stage_1[8][28]), .cin(stage_1[8][29]), .cout(stage_2[9][9]), .s(stage_2[8][23]) );
FA FA_2_129 ( .a(stage_1[8][30]), .b(stage_1[8][31]), .cin(stage_1[8][32]), .cout(stage_2[9][10]), .s(stage_2[8][24]) );
FA FA_2_130 ( .a(stage_1[8][33]), .b(stage_1[8][34]), .cin(stage_1[8][35]), .cout(stage_2[9][11]), .s(stage_2[8][25]) );
FA FA_2_131 ( .a(stage_1[8][36]), .b(stage_1[8][37]), .cin(stage_1[8][38]), .cout(stage_2[9][12]), .s(stage_2[8][26]) );
FA FA_2_132 ( .a(stage_1[8][39]), .b(stage_1[8][40]), .cin(stage_1[8][41]), .cout(stage_2[9][13]), .s(stage_2[8][27]) );
assign stage_2[8][28] = stage_1[8][42];
FA FA_2_133 ( .a(stage_1[9][0]), .b(stage_1[9][1]), .cin(stage_1[9][2]), .cout(stage_2[10][0]), .s(stage_2[9][14]) );
FA FA_2_134 ( .a(stage_1[9][3]), .b(stage_1[9][4]), .cin(stage_1[9][5]), .cout(stage_2[10][1]), .s(stage_2[9][15]) );
FA FA_2_135 ( .a(stage_1[9][6]), .b(stage_1[9][7]), .cin(stage_1[9][8]), .cout(stage_2[10][2]), .s(stage_2[9][16]) );
FA FA_2_136 ( .a(stage_1[9][9]), .b(stage_1[9][10]), .cin(stage_1[9][11]), .cout(stage_2[10][3]), .s(stage_2[9][17]) );
FA FA_2_137 ( .a(stage_1[9][12]), .b(stage_1[9][13]), .cin(stage_1[9][14]), .cout(stage_2[10][4]), .s(stage_2[9][18]) );
FA FA_2_138 ( .a(stage_1[9][15]), .b(stage_1[9][16]), .cin(stage_1[9][17]), .cout(stage_2[10][5]), .s(stage_2[9][19]) );
FA FA_2_139 ( .a(stage_1[9][18]), .b(stage_1[9][19]), .cin(stage_1[9][20]), .cout(stage_2[10][6]), .s(stage_2[9][20]) );
FA FA_2_140 ( .a(stage_1[9][21]), .b(stage_1[9][22]), .cin(stage_1[9][23]), .cout(stage_2[10][7]), .s(stage_2[9][21]) );
FA FA_2_141 ( .a(stage_1[9][24]), .b(stage_1[9][25]), .cin(stage_1[9][26]), .cout(stage_2[10][8]), .s(stage_2[9][22]) );
FA FA_2_142 ( .a(stage_1[9][27]), .b(stage_1[9][28]), .cin(stage_1[9][29]), .cout(stage_2[10][9]), .s(stage_2[9][23]) );
FA FA_2_143 ( .a(stage_1[9][30]), .b(stage_1[9][31]), .cin(stage_1[9][32]), .cout(stage_2[10][10]), .s(stage_2[9][24]) );
FA FA_2_144 ( .a(stage_1[9][33]), .b(stage_1[9][34]), .cin(stage_1[9][35]), .cout(stage_2[10][11]), .s(stage_2[9][25]) );
FA FA_2_145 ( .a(stage_1[9][36]), .b(stage_1[9][37]), .cin(stage_1[9][38]), .cout(stage_2[10][12]), .s(stage_2[9][26]) );
FA FA_2_146 ( .a(stage_1[9][39]), .b(stage_1[9][40]), .cin(stage_1[9][41]), .cout(stage_2[10][13]), .s(stage_2[9][27]) );
assign stage_2[9][28] = stage_1[9][42];
FA FA_2_147 ( .a(stage_1[10][0]), .b(stage_1[10][1]), .cin(stage_1[10][2]), .cout(stage_2[11][0]), .s(stage_2[10][14]) );
FA FA_2_148 ( .a(stage_1[10][3]), .b(stage_1[10][4]), .cin(stage_1[10][5]), .cout(stage_2[11][1]), .s(stage_2[10][15]) );
FA FA_2_149 ( .a(stage_1[10][6]), .b(stage_1[10][7]), .cin(stage_1[10][8]), .cout(stage_2[11][2]), .s(stage_2[10][16]) );
FA FA_2_150 ( .a(stage_1[10][9]), .b(stage_1[10][10]), .cin(stage_1[10][11]), .cout(stage_2[11][3]), .s(stage_2[10][17]) );
FA FA_2_151 ( .a(stage_1[10][12]), .b(stage_1[10][13]), .cin(stage_1[10][14]), .cout(stage_2[11][4]), .s(stage_2[10][18]) );
FA FA_2_152 ( .a(stage_1[10][15]), .b(stage_1[10][16]), .cin(stage_1[10][17]), .cout(stage_2[11][5]), .s(stage_2[10][19]) );
FA FA_2_153 ( .a(stage_1[10][18]), .b(stage_1[10][19]), .cin(stage_1[10][20]), .cout(stage_2[11][6]), .s(stage_2[10][20]) );
FA FA_2_154 ( .a(stage_1[10][21]), .b(stage_1[10][22]), .cin(stage_1[10][23]), .cout(stage_2[11][7]), .s(stage_2[10][21]) );
FA FA_2_155 ( .a(stage_1[10][24]), .b(stage_1[10][25]), .cin(stage_1[10][26]), .cout(stage_2[11][8]), .s(stage_2[10][22]) );
FA FA_2_156 ( .a(stage_1[10][27]), .b(stage_1[10][28]), .cin(stage_1[10][29]), .cout(stage_2[11][9]), .s(stage_2[10][23]) );
FA FA_2_157 ( .a(stage_1[10][30]), .b(stage_1[10][31]), .cin(stage_1[10][32]), .cout(stage_2[11][10]), .s(stage_2[10][24]) );
FA FA_2_158 ( .a(stage_1[10][33]), .b(stage_1[10][34]), .cin(stage_1[10][35]), .cout(stage_2[11][11]), .s(stage_2[10][25]) );
FA FA_2_159 ( .a(stage_1[10][36]), .b(stage_1[10][37]), .cin(stage_1[10][38]), .cout(stage_2[11][12]), .s(stage_2[10][26]) );
FA FA_2_160 ( .a(stage_1[10][39]), .b(stage_1[10][40]), .cin(stage_1[10][41]), .cout(stage_2[11][13]), .s(stage_2[10][27]) );
assign stage_2[10][28] = stage_1[10][42];
FA FA_2_161 ( .a(stage_1[11][0]), .b(stage_1[11][1]), .cin(stage_1[11][2]), .cout(stage_2[12][0]), .s(stage_2[11][14]) );
FA FA_2_162 ( .a(stage_1[11][3]), .b(stage_1[11][4]), .cin(stage_1[11][5]), .cout(stage_2[12][1]), .s(stage_2[11][15]) );
FA FA_2_163 ( .a(stage_1[11][6]), .b(stage_1[11][7]), .cin(stage_1[11][8]), .cout(stage_2[12][2]), .s(stage_2[11][16]) );
FA FA_2_164 ( .a(stage_1[11][9]), .b(stage_1[11][10]), .cin(stage_1[11][11]), .cout(stage_2[12][3]), .s(stage_2[11][17]) );
FA FA_2_165 ( .a(stage_1[11][12]), .b(stage_1[11][13]), .cin(stage_1[11][14]), .cout(stage_2[12][4]), .s(stage_2[11][18]) );
FA FA_2_166 ( .a(stage_1[11][15]), .b(stage_1[11][16]), .cin(stage_1[11][17]), .cout(stage_2[12][5]), .s(stage_2[11][19]) );
FA FA_2_167 ( .a(stage_1[11][18]), .b(stage_1[11][19]), .cin(stage_1[11][20]), .cout(stage_2[12][6]), .s(stage_2[11][20]) );
FA FA_2_168 ( .a(stage_1[11][21]), .b(stage_1[11][22]), .cin(stage_1[11][23]), .cout(stage_2[12][7]), .s(stage_2[11][21]) );
FA FA_2_169 ( .a(stage_1[11][24]), .b(stage_1[11][25]), .cin(stage_1[11][26]), .cout(stage_2[12][8]), .s(stage_2[11][22]) );
FA FA_2_170 ( .a(stage_1[11][27]), .b(stage_1[11][28]), .cin(stage_1[11][29]), .cout(stage_2[12][9]), .s(stage_2[11][23]) );
FA FA_2_171 ( .a(stage_1[11][30]), .b(stage_1[11][31]), .cin(stage_1[11][32]), .cout(stage_2[12][10]), .s(stage_2[11][24]) );
FA FA_2_172 ( .a(stage_1[11][33]), .b(stage_1[11][34]), .cin(stage_1[11][35]), .cout(stage_2[12][11]), .s(stage_2[11][25]) );
FA FA_2_173 ( .a(stage_1[11][36]), .b(stage_1[11][37]), .cin(stage_1[11][38]), .cout(stage_2[12][12]), .s(stage_2[11][26]) );
FA FA_2_174 ( .a(stage_1[11][39]), .b(stage_1[11][40]), .cin(stage_1[11][41]), .cout(stage_2[12][13]), .s(stage_2[11][27]) );
assign stage_2[11][28] = stage_1[11][42];
FA FA_2_175 ( .a(stage_1[12][0]), .b(stage_1[12][1]), .cin(stage_1[12][2]), .cout(stage_2[13][0]), .s(stage_2[12][14]) );
FA FA_2_176 ( .a(stage_1[12][3]), .b(stage_1[12][4]), .cin(stage_1[12][5]), .cout(stage_2[13][1]), .s(stage_2[12][15]) );
FA FA_2_177 ( .a(stage_1[12][6]), .b(stage_1[12][7]), .cin(stage_1[12][8]), .cout(stage_2[13][2]), .s(stage_2[12][16]) );
FA FA_2_178 ( .a(stage_1[12][9]), .b(stage_1[12][10]), .cin(stage_1[12][11]), .cout(stage_2[13][3]), .s(stage_2[12][17]) );
FA FA_2_179 ( .a(stage_1[12][12]), .b(stage_1[12][13]), .cin(stage_1[12][14]), .cout(stage_2[13][4]), .s(stage_2[12][18]) );
FA FA_2_180 ( .a(stage_1[12][15]), .b(stage_1[12][16]), .cin(stage_1[12][17]), .cout(stage_2[13][5]), .s(stage_2[12][19]) );
FA FA_2_181 ( .a(stage_1[12][18]), .b(stage_1[12][19]), .cin(stage_1[12][20]), .cout(stage_2[13][6]), .s(stage_2[12][20]) );
FA FA_2_182 ( .a(stage_1[12][21]), .b(stage_1[12][22]), .cin(stage_1[12][23]), .cout(stage_2[13][7]), .s(stage_2[12][21]) );
FA FA_2_183 ( .a(stage_1[12][24]), .b(stage_1[12][25]), .cin(stage_1[12][26]), .cout(stage_2[13][8]), .s(stage_2[12][22]) );
FA FA_2_184 ( .a(stage_1[12][27]), .b(stage_1[12][28]), .cin(stage_1[12][29]), .cout(stage_2[13][9]), .s(stage_2[12][23]) );
FA FA_2_185 ( .a(stage_1[12][30]), .b(stage_1[12][31]), .cin(stage_1[12][32]), .cout(stage_2[13][10]), .s(stage_2[12][24]) );
FA FA_2_186 ( .a(stage_1[12][33]), .b(stage_1[12][34]), .cin(stage_1[12][35]), .cout(stage_2[13][11]), .s(stage_2[12][25]) );
FA FA_2_187 ( .a(stage_1[12][36]), .b(stage_1[12][37]), .cin(stage_1[12][38]), .cout(stage_2[13][12]), .s(stage_2[12][26]) );
FA FA_2_188 ( .a(stage_1[12][39]), .b(stage_1[12][40]), .cin(stage_1[12][41]), .cout(stage_2[13][13]), .s(stage_2[12][27]) );
assign stage_2[12][28] = stage_1[12][42];
FA FA_2_189 ( .a(stage_1[13][0]), .b(stage_1[13][1]), .cin(stage_1[13][2]), .cout(stage_2[14][0]), .s(stage_2[13][14]) );
FA FA_2_190 ( .a(stage_1[13][3]), .b(stage_1[13][4]), .cin(stage_1[13][5]), .cout(stage_2[14][1]), .s(stage_2[13][15]) );
FA FA_2_191 ( .a(stage_1[13][6]), .b(stage_1[13][7]), .cin(stage_1[13][8]), .cout(stage_2[14][2]), .s(stage_2[13][16]) );
FA FA_2_192 ( .a(stage_1[13][9]), .b(stage_1[13][10]), .cin(stage_1[13][11]), .cout(stage_2[14][3]), .s(stage_2[13][17]) );
FA FA_2_193 ( .a(stage_1[13][12]), .b(stage_1[13][13]), .cin(stage_1[13][14]), .cout(stage_2[14][4]), .s(stage_2[13][18]) );
FA FA_2_194 ( .a(stage_1[13][15]), .b(stage_1[13][16]), .cin(stage_1[13][17]), .cout(stage_2[14][5]), .s(stage_2[13][19]) );
FA FA_2_195 ( .a(stage_1[13][18]), .b(stage_1[13][19]), .cin(stage_1[13][20]), .cout(stage_2[14][6]), .s(stage_2[13][20]) );
FA FA_2_196 ( .a(stage_1[13][21]), .b(stage_1[13][22]), .cin(stage_1[13][23]), .cout(stage_2[14][7]), .s(stage_2[13][21]) );
FA FA_2_197 ( .a(stage_1[13][24]), .b(stage_1[13][25]), .cin(stage_1[13][26]), .cout(stage_2[14][8]), .s(stage_2[13][22]) );
FA FA_2_198 ( .a(stage_1[13][27]), .b(stage_1[13][28]), .cin(stage_1[13][29]), .cout(stage_2[14][9]), .s(stage_2[13][23]) );
FA FA_2_199 ( .a(stage_1[13][30]), .b(stage_1[13][31]), .cin(stage_1[13][32]), .cout(stage_2[14][10]), .s(stage_2[13][24]) );
FA FA_2_200 ( .a(stage_1[13][33]), .b(stage_1[13][34]), .cin(stage_1[13][35]), .cout(stage_2[14][11]), .s(stage_2[13][25]) );
FA FA_2_201 ( .a(stage_1[13][36]), .b(stage_1[13][37]), .cin(stage_1[13][38]), .cout(stage_2[14][12]), .s(stage_2[13][26]) );
FA FA_2_202 ( .a(stage_1[13][39]), .b(stage_1[13][40]), .cin(stage_1[13][41]), .cout(stage_2[14][13]), .s(stage_2[13][27]) );
assign stage_2[13][28] = stage_1[13][42];
FA FA_2_203 ( .a(stage_1[14][0]), .b(stage_1[14][1]), .cin(stage_1[14][2]), .cout(stage_2[15][0]), .s(stage_2[14][14]) );
FA FA_2_204 ( .a(stage_1[14][3]), .b(stage_1[14][4]), .cin(stage_1[14][5]), .cout(stage_2[15][1]), .s(stage_2[14][15]) );
FA FA_2_205 ( .a(stage_1[14][6]), .b(stage_1[14][7]), .cin(stage_1[14][8]), .cout(stage_2[15][2]), .s(stage_2[14][16]) );
FA FA_2_206 ( .a(stage_1[14][9]), .b(stage_1[14][10]), .cin(stage_1[14][11]), .cout(stage_2[15][3]), .s(stage_2[14][17]) );
FA FA_2_207 ( .a(stage_1[14][12]), .b(stage_1[14][13]), .cin(stage_1[14][14]), .cout(stage_2[15][4]), .s(stage_2[14][18]) );
FA FA_2_208 ( .a(stage_1[14][15]), .b(stage_1[14][16]), .cin(stage_1[14][17]), .cout(stage_2[15][5]), .s(stage_2[14][19]) );
FA FA_2_209 ( .a(stage_1[14][18]), .b(stage_1[14][19]), .cin(stage_1[14][20]), .cout(stage_2[15][6]), .s(stage_2[14][20]) );
FA FA_2_210 ( .a(stage_1[14][21]), .b(stage_1[14][22]), .cin(stage_1[14][23]), .cout(stage_2[15][7]), .s(stage_2[14][21]) );
FA FA_2_211 ( .a(stage_1[14][24]), .b(stage_1[14][25]), .cin(stage_1[14][26]), .cout(stage_2[15][8]), .s(stage_2[14][22]) );
FA FA_2_212 ( .a(stage_1[14][27]), .b(stage_1[14][28]), .cin(stage_1[14][29]), .cout(stage_2[15][9]), .s(stage_2[14][23]) );
FA FA_2_213 ( .a(stage_1[14][30]), .b(stage_1[14][31]), .cin(stage_1[14][32]), .cout(stage_2[15][10]), .s(stage_2[14][24]) );
FA FA_2_214 ( .a(stage_1[14][33]), .b(stage_1[14][34]), .cin(stage_1[14][35]), .cout(stage_2[15][11]), .s(stage_2[14][25]) );
FA FA_2_215 ( .a(stage_1[14][36]), .b(stage_1[14][37]), .cin(stage_1[14][38]), .cout(stage_2[15][12]), .s(stage_2[14][26]) );
FA FA_2_216 ( .a(stage_1[14][39]), .b(stage_1[14][40]), .cin(stage_1[14][41]), .cout(stage_2[15][13]), .s(stage_2[14][27]) );
assign stage_2[14][28] = stage_1[14][42];
FA FA_2_217 ( .a(stage_1[15][0]), .b(stage_1[15][1]), .cin(stage_1[15][2]), .cout(stage_2[16][0]), .s(stage_2[15][14]) );
FA FA_2_218 ( .a(stage_1[15][3]), .b(stage_1[15][4]), .cin(stage_1[15][5]), .cout(stage_2[16][1]), .s(stage_2[15][15]) );
FA FA_2_219 ( .a(stage_1[15][6]), .b(stage_1[15][7]), .cin(stage_1[15][8]), .cout(stage_2[16][2]), .s(stage_2[15][16]) );
FA FA_2_220 ( .a(stage_1[15][9]), .b(stage_1[15][10]), .cin(stage_1[15][11]), .cout(stage_2[16][3]), .s(stage_2[15][17]) );
FA FA_2_221 ( .a(stage_1[15][12]), .b(stage_1[15][13]), .cin(stage_1[15][14]), .cout(stage_2[16][4]), .s(stage_2[15][18]) );
FA FA_2_222 ( .a(stage_1[15][15]), .b(stage_1[15][16]), .cin(stage_1[15][17]), .cout(stage_2[16][5]), .s(stage_2[15][19]) );
FA FA_2_223 ( .a(stage_1[15][18]), .b(stage_1[15][19]), .cin(stage_1[15][20]), .cout(stage_2[16][6]), .s(stage_2[15][20]) );
FA FA_2_224 ( .a(stage_1[15][21]), .b(stage_1[15][22]), .cin(stage_1[15][23]), .cout(stage_2[16][7]), .s(stage_2[15][21]) );
FA FA_2_225 ( .a(stage_1[15][24]), .b(stage_1[15][25]), .cin(stage_1[15][26]), .cout(stage_2[16][8]), .s(stage_2[15][22]) );
FA FA_2_226 ( .a(stage_1[15][27]), .b(stage_1[15][28]), .cin(stage_1[15][29]), .cout(stage_2[16][9]), .s(stage_2[15][23]) );
FA FA_2_227 ( .a(stage_1[15][30]), .b(stage_1[15][31]), .cin(stage_1[15][32]), .cout(stage_2[16][10]), .s(stage_2[15][24]) );
FA FA_2_228 ( .a(stage_1[15][33]), .b(stage_1[15][34]), .cin(stage_1[15][35]), .cout(stage_2[16][11]), .s(stage_2[15][25]) );
FA FA_2_229 ( .a(stage_1[15][36]), .b(stage_1[15][37]), .cin(stage_1[15][38]), .cout(stage_2[16][12]), .s(stage_2[15][26]) );
FA FA_2_230 ( .a(stage_1[15][39]), .b(stage_1[15][40]), .cin(stage_1[15][41]), .cout(stage_2[16][13]), .s(stage_2[15][27]) );
assign stage_2[15][28] = stage_1[15][42];
FA FA_2_231 ( .a(stage_1[16][0]), .b(stage_1[16][1]), .cin(stage_1[16][2]), .cout(stage_2[17][0]), .s(stage_2[16][14]) );
FA FA_2_232 ( .a(stage_1[16][3]), .b(stage_1[16][4]), .cin(stage_1[16][5]), .cout(stage_2[17][1]), .s(stage_2[16][15]) );
FA FA_2_233 ( .a(stage_1[16][6]), .b(stage_1[16][7]), .cin(stage_1[16][8]), .cout(stage_2[17][2]), .s(stage_2[16][16]) );
FA FA_2_234 ( .a(stage_1[16][9]), .b(stage_1[16][10]), .cin(stage_1[16][11]), .cout(stage_2[17][3]), .s(stage_2[16][17]) );
FA FA_2_235 ( .a(stage_1[16][12]), .b(stage_1[16][13]), .cin(stage_1[16][14]), .cout(stage_2[17][4]), .s(stage_2[16][18]) );
FA FA_2_236 ( .a(stage_1[16][15]), .b(stage_1[16][16]), .cin(stage_1[16][17]), .cout(stage_2[17][5]), .s(stage_2[16][19]) );
FA FA_2_237 ( .a(stage_1[16][18]), .b(stage_1[16][19]), .cin(stage_1[16][20]), .cout(stage_2[17][6]), .s(stage_2[16][20]) );

wire stage_3 [`NBIT+3:0][`NDATA*2:0];
FA FA_3_0 ( .a(stage_2[0][0]), .b(stage_2[0][1]), .cin(stage_2[0][2]), .cout(stage_3[1][0]), .s(stage_3[0][0]) );
FA FA_3_1 ( .a(stage_2[0][3]), .b(stage_2[0][4]), .cin(stage_2[0][5]), .cout(stage_3[1][1]), .s(stage_3[0][1]) );
FA FA_3_2 ( .a(stage_2[0][6]), .b(stage_2[0][7]), .cin(stage_2[0][8]), .cout(stage_3[1][2]), .s(stage_3[0][2]) );
FA FA_3_3 ( .a(stage_2[0][9]), .b(stage_2[0][10]), .cin(stage_2[0][11]), .cout(stage_3[1][3]), .s(stage_3[0][3]) );
FA FA_3_4 ( .a(stage_2[0][12]), .b(stage_2[0][13]), .cin(stage_2[0][14]), .cout(stage_3[1][4]), .s(stage_3[0][4]) );
FA FA_3_5 ( .a(stage_2[1][0]), .b(stage_2[1][1]), .cin(stage_2[1][2]), .cout(stage_3[2][0]), .s(stage_3[1][5]) );
FA FA_3_6 ( .a(stage_2[1][3]), .b(stage_2[1][4]), .cin(stage_2[1][5]), .cout(stage_3[2][1]), .s(stage_3[1][6]) );
FA FA_3_7 ( .a(stage_2[1][6]), .b(stage_2[1][7]), .cin(stage_2[1][8]), .cout(stage_3[2][2]), .s(stage_3[1][7]) );
FA FA_3_8 ( .a(stage_2[1][9]), .b(stage_2[1][10]), .cin(stage_2[1][11]), .cout(stage_3[2][3]), .s(stage_3[1][8]) );
FA FA_3_9 ( .a(stage_2[1][12]), .b(stage_2[1][13]), .cin(stage_2[1][14]), .cout(stage_3[2][4]), .s(stage_3[1][9]) );
FA FA_3_10 ( .a(stage_2[1][15]), .b(stage_2[1][16]), .cin(stage_2[1][17]), .cout(stage_3[2][5]), .s(stage_3[1][10]) );
FA FA_3_11 ( .a(stage_2[1][18]), .b(stage_2[1][19]), .cin(stage_2[1][20]), .cout(stage_3[2][6]), .s(stage_3[1][11]) );
FA FA_3_12 ( .a(stage_2[1][21]), .b(stage_2[1][22]), .cin(stage_2[1][23]), .cout(stage_3[2][7]), .s(stage_3[1][12]) );
FA FA_3_13 ( .a(stage_2[1][24]), .b(stage_2[1][25]), .cin(stage_2[1][26]), .cout(stage_3[2][8]), .s(stage_3[1][13]) );
FA FA_3_14 ( .a(stage_2[1][27]), .b(stage_2[1][28]), .cin(stage_2[1][29]), .cout(stage_3[2][9]), .s(stage_3[1][14]) );
FA FA_3_15 ( .a(stage_2[1][30]), .b(stage_2[1][31]), .cin(stage_2[1][32]), .cout(stage_3[2][10]), .s(stage_3[1][15]) );
FA FA_3_16 ( .a(stage_2[1][33]), .b(stage_2[1][34]), .cin(stage_2[1][35]), .cout(stage_3[2][11]), .s(stage_3[1][16]) );
FA FA_3_17 ( .a(stage_2[2][0]), .b(stage_2[2][1]), .cin(stage_2[2][2]), .cout(stage_3[3][0]), .s(stage_3[2][12]) );
FA FA_3_18 ( .a(stage_2[2][3]), .b(stage_2[2][4]), .cin(stage_2[2][5]), .cout(stage_3[3][1]), .s(stage_3[2][13]) );
FA FA_3_19 ( .a(stage_2[2][6]), .b(stage_2[2][7]), .cin(stage_2[2][8]), .cout(stage_3[3][2]), .s(stage_3[2][14]) );
FA FA_3_20 ( .a(stage_2[2][9]), .b(stage_2[2][10]), .cin(stage_2[2][11]), .cout(stage_3[3][3]), .s(stage_3[2][15]) );
FA FA_3_21 ( .a(stage_2[2][12]), .b(stage_2[2][13]), .cin(stage_2[2][14]), .cout(stage_3[3][4]), .s(stage_3[2][16]) );
FA FA_3_22 ( .a(stage_2[2][15]), .b(stage_2[2][16]), .cin(stage_2[2][17]), .cout(stage_3[3][5]), .s(stage_3[2][17]) );
FA FA_3_23 ( .a(stage_2[2][18]), .b(stage_2[2][19]), .cin(stage_2[2][20]), .cout(stage_3[3][6]), .s(stage_3[2][18]) );
FA FA_3_24 ( .a(stage_2[2][21]), .b(stage_2[2][22]), .cin(stage_2[2][23]), .cout(stage_3[3][7]), .s(stage_3[2][19]) );
FA FA_3_25 ( .a(stage_2[2][24]), .b(stage_2[2][25]), .cin(stage_2[2][26]), .cout(stage_3[3][8]), .s(stage_3[2][20]) );
FA FA_3_26 ( .a(stage_2[2][27]), .b(stage_2[2][28]), .cin(stage_2[2][29]), .cout(stage_3[3][9]), .s(stage_3[2][21]) );
FA FA_3_27 ( .a(stage_2[2][30]), .b(stage_2[2][31]), .cin(stage_2[2][32]), .cout(stage_3[3][10]), .s(stage_3[2][22]) );
FA FA_3_28 ( .a(stage_2[2][33]), .b(stage_2[2][34]), .cin(stage_2[2][35]), .cout(stage_3[3][11]), .s(stage_3[2][23]) );
assign stage_3[2][24] = stage_2[2][36];
FA FA_3_29 ( .a(stage_2[3][0]), .b(stage_2[3][1]), .cin(stage_2[3][2]), .cout(stage_3[4][0]), .s(stage_3[3][12]) );
FA FA_3_30 ( .a(stage_2[3][3]), .b(stage_2[3][4]), .cin(stage_2[3][5]), .cout(stage_3[4][1]), .s(stage_3[3][13]) );
FA FA_3_31 ( .a(stage_2[3][6]), .b(stage_2[3][7]), .cin(stage_2[3][8]), .cout(stage_3[4][2]), .s(stage_3[3][14]) );
FA FA_3_32 ( .a(stage_2[3][9]), .b(stage_2[3][10]), .cin(stage_2[3][11]), .cout(stage_3[4][3]), .s(stage_3[3][15]) );
FA FA_3_33 ( .a(stage_2[3][12]), .b(stage_2[3][13]), .cin(stage_2[3][14]), .cout(stage_3[4][4]), .s(stage_3[3][16]) );
FA FA_3_34 ( .a(stage_2[3][15]), .b(stage_2[3][16]), .cin(stage_2[3][17]), .cout(stage_3[4][5]), .s(stage_3[3][17]) );
FA FA_3_35 ( .a(stage_2[3][18]), .b(stage_2[3][19]), .cin(stage_2[3][20]), .cout(stage_3[4][6]), .s(stage_3[3][18]) );
FA FA_3_36 ( .a(stage_2[3][21]), .b(stage_2[3][22]), .cin(stage_2[3][23]), .cout(stage_3[4][7]), .s(stage_3[3][19]) );
FA FA_3_37 ( .a(stage_2[3][24]), .b(stage_2[3][25]), .cin(stage_2[3][26]), .cout(stage_3[4][8]), .s(stage_3[3][20]) );
HA HA_3_0 ( .a(stage_2[3][27]), .b(stage_2[3][28]), .cout(stage_3[4][9]), .s(stage_3[3][21]) );
FA FA_3_38 ( .a(stage_2[4][0]), .b(stage_2[4][1]), .cin(stage_2[4][2]), .cout(stage_3[5][0]), .s(stage_3[4][10]) );
FA FA_3_39 ( .a(stage_2[4][3]), .b(stage_2[4][4]), .cin(stage_2[4][5]), .cout(stage_3[5][1]), .s(stage_3[4][11]) );
FA FA_3_40 ( .a(stage_2[4][6]), .b(stage_2[4][7]), .cin(stage_2[4][8]), .cout(stage_3[5][2]), .s(stage_3[4][12]) );
FA FA_3_41 ( .a(stage_2[4][9]), .b(stage_2[4][10]), .cin(stage_2[4][11]), .cout(stage_3[5][3]), .s(stage_3[4][13]) );
FA FA_3_42 ( .a(stage_2[4][12]), .b(stage_2[4][13]), .cin(stage_2[4][14]), .cout(stage_3[5][4]), .s(stage_3[4][14]) );
FA FA_3_43 ( .a(stage_2[4][15]), .b(stage_2[4][16]), .cin(stage_2[4][17]), .cout(stage_3[5][5]), .s(stage_3[4][15]) );
FA FA_3_44 ( .a(stage_2[4][18]), .b(stage_2[4][19]), .cin(stage_2[4][20]), .cout(stage_3[5][6]), .s(stage_3[4][16]) );
FA FA_3_45 ( .a(stage_2[4][21]), .b(stage_2[4][22]), .cin(stage_2[4][23]), .cout(stage_3[5][7]), .s(stage_3[4][17]) );
FA FA_3_46 ( .a(stage_2[4][24]), .b(stage_2[4][25]), .cin(stage_2[4][26]), .cout(stage_3[5][8]), .s(stage_3[4][18]) );
HA HA_3_1 ( .a(stage_2[4][27]), .b(stage_2[4][28]), .cout(stage_3[5][9]), .s(stage_3[4][19]) );
FA FA_3_47 ( .a(stage_2[5][0]), .b(stage_2[5][1]), .cin(stage_2[5][2]), .cout(stage_3[6][0]), .s(stage_3[5][10]) );
FA FA_3_48 ( .a(stage_2[5][3]), .b(stage_2[5][4]), .cin(stage_2[5][5]), .cout(stage_3[6][1]), .s(stage_3[5][11]) );
FA FA_3_49 ( .a(stage_2[5][6]), .b(stage_2[5][7]), .cin(stage_2[5][8]), .cout(stage_3[6][2]), .s(stage_3[5][12]) );
FA FA_3_50 ( .a(stage_2[5][9]), .b(stage_2[5][10]), .cin(stage_2[5][11]), .cout(stage_3[6][3]), .s(stage_3[5][13]) );
FA FA_3_51 ( .a(stage_2[5][12]), .b(stage_2[5][13]), .cin(stage_2[5][14]), .cout(stage_3[6][4]), .s(stage_3[5][14]) );
FA FA_3_52 ( .a(stage_2[5][15]), .b(stage_2[5][16]), .cin(stage_2[5][17]), .cout(stage_3[6][5]), .s(stage_3[5][15]) );
FA FA_3_53 ( .a(stage_2[5][18]), .b(stage_2[5][19]), .cin(stage_2[5][20]), .cout(stage_3[6][6]), .s(stage_3[5][16]) );
FA FA_3_54 ( .a(stage_2[5][21]), .b(stage_2[5][22]), .cin(stage_2[5][23]), .cout(stage_3[6][7]), .s(stage_3[5][17]) );
FA FA_3_55 ( .a(stage_2[5][24]), .b(stage_2[5][25]), .cin(stage_2[5][26]), .cout(stage_3[6][8]), .s(stage_3[5][18]) );
HA HA_3_2 ( .a(stage_2[5][27]), .b(stage_2[5][28]), .cout(stage_3[6][9]), .s(stage_3[5][19]) );
FA FA_3_56 ( .a(stage_2[6][0]), .b(stage_2[6][1]), .cin(stage_2[6][2]), .cout(stage_3[7][0]), .s(stage_3[6][10]) );
FA FA_3_57 ( .a(stage_2[6][3]), .b(stage_2[6][4]), .cin(stage_2[6][5]), .cout(stage_3[7][1]), .s(stage_3[6][11]) );
FA FA_3_58 ( .a(stage_2[6][6]), .b(stage_2[6][7]), .cin(stage_2[6][8]), .cout(stage_3[7][2]), .s(stage_3[6][12]) );
FA FA_3_59 ( .a(stage_2[6][9]), .b(stage_2[6][10]), .cin(stage_2[6][11]), .cout(stage_3[7][3]), .s(stage_3[6][13]) );
FA FA_3_60 ( .a(stage_2[6][12]), .b(stage_2[6][13]), .cin(stage_2[6][14]), .cout(stage_3[7][4]), .s(stage_3[6][14]) );
FA FA_3_61 ( .a(stage_2[6][15]), .b(stage_2[6][16]), .cin(stage_2[6][17]), .cout(stage_3[7][5]), .s(stage_3[6][15]) );
FA FA_3_62 ( .a(stage_2[6][18]), .b(stage_2[6][19]), .cin(stage_2[6][20]), .cout(stage_3[7][6]), .s(stage_3[6][16]) );
FA FA_3_63 ( .a(stage_2[6][21]), .b(stage_2[6][22]), .cin(stage_2[6][23]), .cout(stage_3[7][7]), .s(stage_3[6][17]) );
FA FA_3_64 ( .a(stage_2[6][24]), .b(stage_2[6][25]), .cin(stage_2[6][26]), .cout(stage_3[7][8]), .s(stage_3[6][18]) );
HA HA_3_3 ( .a(stage_2[6][27]), .b(stage_2[6][28]), .cout(stage_3[7][9]), .s(stage_3[6][19]) );
FA FA_3_65 ( .a(stage_2[7][0]), .b(stage_2[7][1]), .cin(stage_2[7][2]), .cout(stage_3[8][0]), .s(stage_3[7][10]) );
FA FA_3_66 ( .a(stage_2[7][3]), .b(stage_2[7][4]), .cin(stage_2[7][5]), .cout(stage_3[8][1]), .s(stage_3[7][11]) );
FA FA_3_67 ( .a(stage_2[7][6]), .b(stage_2[7][7]), .cin(stage_2[7][8]), .cout(stage_3[8][2]), .s(stage_3[7][12]) );
FA FA_3_68 ( .a(stage_2[7][9]), .b(stage_2[7][10]), .cin(stage_2[7][11]), .cout(stage_3[8][3]), .s(stage_3[7][13]) );
FA FA_3_69 ( .a(stage_2[7][12]), .b(stage_2[7][13]), .cin(stage_2[7][14]), .cout(stage_3[8][4]), .s(stage_3[7][14]) );
FA FA_3_70 ( .a(stage_2[7][15]), .b(stage_2[7][16]), .cin(stage_2[7][17]), .cout(stage_3[8][5]), .s(stage_3[7][15]) );
FA FA_3_71 ( .a(stage_2[7][18]), .b(stage_2[7][19]), .cin(stage_2[7][20]), .cout(stage_3[8][6]), .s(stage_3[7][16]) );
FA FA_3_72 ( .a(stage_2[7][21]), .b(stage_2[7][22]), .cin(stage_2[7][23]), .cout(stage_3[8][7]), .s(stage_3[7][17]) );
FA FA_3_73 ( .a(stage_2[7][24]), .b(stage_2[7][25]), .cin(stage_2[7][26]), .cout(stage_3[8][8]), .s(stage_3[7][18]) );
HA HA_3_4 ( .a(stage_2[7][27]), .b(stage_2[7][28]), .cout(stage_3[8][9]), .s(stage_3[7][19]) );
FA FA_3_74 ( .a(stage_2[8][0]), .b(stage_2[8][1]), .cin(stage_2[8][2]), .cout(stage_3[9][0]), .s(stage_3[8][10]) );
FA FA_3_75 ( .a(stage_2[8][3]), .b(stage_2[8][4]), .cin(stage_2[8][5]), .cout(stage_3[9][1]), .s(stage_3[8][11]) );
FA FA_3_76 ( .a(stage_2[8][6]), .b(stage_2[8][7]), .cin(stage_2[8][8]), .cout(stage_3[9][2]), .s(stage_3[8][12]) );
FA FA_3_77 ( .a(stage_2[8][9]), .b(stage_2[8][10]), .cin(stage_2[8][11]), .cout(stage_3[9][3]), .s(stage_3[8][13]) );
FA FA_3_78 ( .a(stage_2[8][12]), .b(stage_2[8][13]), .cin(stage_2[8][14]), .cout(stage_3[9][4]), .s(stage_3[8][14]) );
FA FA_3_79 ( .a(stage_2[8][15]), .b(stage_2[8][16]), .cin(stage_2[8][17]), .cout(stage_3[9][5]), .s(stage_3[8][15]) );
FA FA_3_80 ( .a(stage_2[8][18]), .b(stage_2[8][19]), .cin(stage_2[8][20]), .cout(stage_3[9][6]), .s(stage_3[8][16]) );
FA FA_3_81 ( .a(stage_2[8][21]), .b(stage_2[8][22]), .cin(stage_2[8][23]), .cout(stage_3[9][7]), .s(stage_3[8][17]) );
FA FA_3_82 ( .a(stage_2[8][24]), .b(stage_2[8][25]), .cin(stage_2[8][26]), .cout(stage_3[9][8]), .s(stage_3[8][18]) );
HA HA_3_5 ( .a(stage_2[8][27]), .b(stage_2[8][28]), .cout(stage_3[9][9]), .s(stage_3[8][19]) );
FA FA_3_83 ( .a(stage_2[9][0]), .b(stage_2[9][1]), .cin(stage_2[9][2]), .cout(stage_3[10][0]), .s(stage_3[9][10]) );
FA FA_3_84 ( .a(stage_2[9][3]), .b(stage_2[9][4]), .cin(stage_2[9][5]), .cout(stage_3[10][1]), .s(stage_3[9][11]) );
FA FA_3_85 ( .a(stage_2[9][6]), .b(stage_2[9][7]), .cin(stage_2[9][8]), .cout(stage_3[10][2]), .s(stage_3[9][12]) );
FA FA_3_86 ( .a(stage_2[9][9]), .b(stage_2[9][10]), .cin(stage_2[9][11]), .cout(stage_3[10][3]), .s(stage_3[9][13]) );
FA FA_3_87 ( .a(stage_2[9][12]), .b(stage_2[9][13]), .cin(stage_2[9][14]), .cout(stage_3[10][4]), .s(stage_3[9][14]) );
FA FA_3_88 ( .a(stage_2[9][15]), .b(stage_2[9][16]), .cin(stage_2[9][17]), .cout(stage_3[10][5]), .s(stage_3[9][15]) );
FA FA_3_89 ( .a(stage_2[9][18]), .b(stage_2[9][19]), .cin(stage_2[9][20]), .cout(stage_3[10][6]), .s(stage_3[9][16]) );
FA FA_3_90 ( .a(stage_2[9][21]), .b(stage_2[9][22]), .cin(stage_2[9][23]), .cout(stage_3[10][7]), .s(stage_3[9][17]) );
FA FA_3_91 ( .a(stage_2[9][24]), .b(stage_2[9][25]), .cin(stage_2[9][26]), .cout(stage_3[10][8]), .s(stage_3[9][18]) );
HA HA_3_6 ( .a(stage_2[9][27]), .b(stage_2[9][28]), .cout(stage_3[10][9]), .s(stage_3[9][19]) );
FA FA_3_92 ( .a(stage_2[10][0]), .b(stage_2[10][1]), .cin(stage_2[10][2]), .cout(stage_3[11][0]), .s(stage_3[10][10]) );
FA FA_3_93 ( .a(stage_2[10][3]), .b(stage_2[10][4]), .cin(stage_2[10][5]), .cout(stage_3[11][1]), .s(stage_3[10][11]) );
FA FA_3_94 ( .a(stage_2[10][6]), .b(stage_2[10][7]), .cin(stage_2[10][8]), .cout(stage_3[11][2]), .s(stage_3[10][12]) );
FA FA_3_95 ( .a(stage_2[10][9]), .b(stage_2[10][10]), .cin(stage_2[10][11]), .cout(stage_3[11][3]), .s(stage_3[10][13]) );
FA FA_3_96 ( .a(stage_2[10][12]), .b(stage_2[10][13]), .cin(stage_2[10][14]), .cout(stage_3[11][4]), .s(stage_3[10][14]) );
FA FA_3_97 ( .a(stage_2[10][15]), .b(stage_2[10][16]), .cin(stage_2[10][17]), .cout(stage_3[11][5]), .s(stage_3[10][15]) );
FA FA_3_98 ( .a(stage_2[10][18]), .b(stage_2[10][19]), .cin(stage_2[10][20]), .cout(stage_3[11][6]), .s(stage_3[10][16]) );
FA FA_3_99 ( .a(stage_2[10][21]), .b(stage_2[10][22]), .cin(stage_2[10][23]), .cout(stage_3[11][7]), .s(stage_3[10][17]) );
FA FA_3_100 ( .a(stage_2[10][24]), .b(stage_2[10][25]), .cin(stage_2[10][26]), .cout(stage_3[11][8]), .s(stage_3[10][18]) );
HA HA_3_7 ( .a(stage_2[10][27]), .b(stage_2[10][28]), .cout(stage_3[11][9]), .s(stage_3[10][19]) );
FA FA_3_101 ( .a(stage_2[11][0]), .b(stage_2[11][1]), .cin(stage_2[11][2]), .cout(stage_3[12][0]), .s(stage_3[11][10]) );
FA FA_3_102 ( .a(stage_2[11][3]), .b(stage_2[11][4]), .cin(stage_2[11][5]), .cout(stage_3[12][1]), .s(stage_3[11][11]) );
FA FA_3_103 ( .a(stage_2[11][6]), .b(stage_2[11][7]), .cin(stage_2[11][8]), .cout(stage_3[12][2]), .s(stage_3[11][12]) );
FA FA_3_104 ( .a(stage_2[11][9]), .b(stage_2[11][10]), .cin(stage_2[11][11]), .cout(stage_3[12][3]), .s(stage_3[11][13]) );
FA FA_3_105 ( .a(stage_2[11][12]), .b(stage_2[11][13]), .cin(stage_2[11][14]), .cout(stage_3[12][4]), .s(stage_3[11][14]) );
FA FA_3_106 ( .a(stage_2[11][15]), .b(stage_2[11][16]), .cin(stage_2[11][17]), .cout(stage_3[12][5]), .s(stage_3[11][15]) );
FA FA_3_107 ( .a(stage_2[11][18]), .b(stage_2[11][19]), .cin(stage_2[11][20]), .cout(stage_3[12][6]), .s(stage_3[11][16]) );
FA FA_3_108 ( .a(stage_2[11][21]), .b(stage_2[11][22]), .cin(stage_2[11][23]), .cout(stage_3[12][7]), .s(stage_3[11][17]) );
FA FA_3_109 ( .a(stage_2[11][24]), .b(stage_2[11][25]), .cin(stage_2[11][26]), .cout(stage_3[12][8]), .s(stage_3[11][18]) );
HA HA_3_8 ( .a(stage_2[11][27]), .b(stage_2[11][28]), .cout(stage_3[12][9]), .s(stage_3[11][19]) );
FA FA_3_110 ( .a(stage_2[12][0]), .b(stage_2[12][1]), .cin(stage_2[12][2]), .cout(stage_3[13][0]), .s(stage_3[12][10]) );
FA FA_3_111 ( .a(stage_2[12][3]), .b(stage_2[12][4]), .cin(stage_2[12][5]), .cout(stage_3[13][1]), .s(stage_3[12][11]) );
FA FA_3_112 ( .a(stage_2[12][6]), .b(stage_2[12][7]), .cin(stage_2[12][8]), .cout(stage_3[13][2]), .s(stage_3[12][12]) );
FA FA_3_113 ( .a(stage_2[12][9]), .b(stage_2[12][10]), .cin(stage_2[12][11]), .cout(stage_3[13][3]), .s(stage_3[12][13]) );
FA FA_3_114 ( .a(stage_2[12][12]), .b(stage_2[12][13]), .cin(stage_2[12][14]), .cout(stage_3[13][4]), .s(stage_3[12][14]) );
FA FA_3_115 ( .a(stage_2[12][15]), .b(stage_2[12][16]), .cin(stage_2[12][17]), .cout(stage_3[13][5]), .s(stage_3[12][15]) );
FA FA_3_116 ( .a(stage_2[12][18]), .b(stage_2[12][19]), .cin(stage_2[12][20]), .cout(stage_3[13][6]), .s(stage_3[12][16]) );
FA FA_3_117 ( .a(stage_2[12][21]), .b(stage_2[12][22]), .cin(stage_2[12][23]), .cout(stage_3[13][7]), .s(stage_3[12][17]) );
FA FA_3_118 ( .a(stage_2[12][24]), .b(stage_2[12][25]), .cin(stage_2[12][26]), .cout(stage_3[13][8]), .s(stage_3[12][18]) );
HA HA_3_9 ( .a(stage_2[12][27]), .b(stage_2[12][28]), .cout(stage_3[13][9]), .s(stage_3[12][19]) );
FA FA_3_119 ( .a(stage_2[13][0]), .b(stage_2[13][1]), .cin(stage_2[13][2]), .cout(stage_3[14][0]), .s(stage_3[13][10]) );
FA FA_3_120 ( .a(stage_2[13][3]), .b(stage_2[13][4]), .cin(stage_2[13][5]), .cout(stage_3[14][1]), .s(stage_3[13][11]) );
FA FA_3_121 ( .a(stage_2[13][6]), .b(stage_2[13][7]), .cin(stage_2[13][8]), .cout(stage_3[14][2]), .s(stage_3[13][12]) );
FA FA_3_122 ( .a(stage_2[13][9]), .b(stage_2[13][10]), .cin(stage_2[13][11]), .cout(stage_3[14][3]), .s(stage_3[13][13]) );
FA FA_3_123 ( .a(stage_2[13][12]), .b(stage_2[13][13]), .cin(stage_2[13][14]), .cout(stage_3[14][4]), .s(stage_3[13][14]) );
FA FA_3_124 ( .a(stage_2[13][15]), .b(stage_2[13][16]), .cin(stage_2[13][17]), .cout(stage_3[14][5]), .s(stage_3[13][15]) );
FA FA_3_125 ( .a(stage_2[13][18]), .b(stage_2[13][19]), .cin(stage_2[13][20]), .cout(stage_3[14][6]), .s(stage_3[13][16]) );
FA FA_3_126 ( .a(stage_2[13][21]), .b(stage_2[13][22]), .cin(stage_2[13][23]), .cout(stage_3[14][7]), .s(stage_3[13][17]) );
FA FA_3_127 ( .a(stage_2[13][24]), .b(stage_2[13][25]), .cin(stage_2[13][26]), .cout(stage_3[14][8]), .s(stage_3[13][18]) );
HA HA_3_10 ( .a(stage_2[13][27]), .b(stage_2[13][28]), .cout(stage_3[14][9]), .s(stage_3[13][19]) );
FA FA_3_128 ( .a(stage_2[14][0]), .b(stage_2[14][1]), .cin(stage_2[14][2]), .cout(stage_3[15][0]), .s(stage_3[14][10]) );
FA FA_3_129 ( .a(stage_2[14][3]), .b(stage_2[14][4]), .cin(stage_2[14][5]), .cout(stage_3[15][1]), .s(stage_3[14][11]) );
FA FA_3_130 ( .a(stage_2[14][6]), .b(stage_2[14][7]), .cin(stage_2[14][8]), .cout(stage_3[15][2]), .s(stage_3[14][12]) );
FA FA_3_131 ( .a(stage_2[14][9]), .b(stage_2[14][10]), .cin(stage_2[14][11]), .cout(stage_3[15][3]), .s(stage_3[14][13]) );
FA FA_3_132 ( .a(stage_2[14][12]), .b(stage_2[14][13]), .cin(stage_2[14][14]), .cout(stage_3[15][4]), .s(stage_3[14][14]) );
FA FA_3_133 ( .a(stage_2[14][15]), .b(stage_2[14][16]), .cin(stage_2[14][17]), .cout(stage_3[15][5]), .s(stage_3[14][15]) );
FA FA_3_134 ( .a(stage_2[14][18]), .b(stage_2[14][19]), .cin(stage_2[14][20]), .cout(stage_3[15][6]), .s(stage_3[14][16]) );
FA FA_3_135 ( .a(stage_2[14][21]), .b(stage_2[14][22]), .cin(stage_2[14][23]), .cout(stage_3[15][7]), .s(stage_3[14][17]) );
FA FA_3_136 ( .a(stage_2[14][24]), .b(stage_2[14][25]), .cin(stage_2[14][26]), .cout(stage_3[15][8]), .s(stage_3[14][18]) );
HA HA_3_11 ( .a(stage_2[14][27]), .b(stage_2[14][28]), .cout(stage_3[15][9]), .s(stage_3[14][19]) );
FA FA_3_137 ( .a(stage_2[15][0]), .b(stage_2[15][1]), .cin(stage_2[15][2]), .cout(stage_3[16][0]), .s(stage_3[15][10]) );
FA FA_3_138 ( .a(stage_2[15][3]), .b(stage_2[15][4]), .cin(stage_2[15][5]), .cout(stage_3[16][1]), .s(stage_3[15][11]) );
FA FA_3_139 ( .a(stage_2[15][6]), .b(stage_2[15][7]), .cin(stage_2[15][8]), .cout(stage_3[16][2]), .s(stage_3[15][12]) );
FA FA_3_140 ( .a(stage_2[15][9]), .b(stage_2[15][10]), .cin(stage_2[15][11]), .cout(stage_3[16][3]), .s(stage_3[15][13]) );
FA FA_3_141 ( .a(stage_2[15][12]), .b(stage_2[15][13]), .cin(stage_2[15][14]), .cout(stage_3[16][4]), .s(stage_3[15][14]) );
FA FA_3_142 ( .a(stage_2[15][15]), .b(stage_2[15][16]), .cin(stage_2[15][17]), .cout(stage_3[16][5]), .s(stage_3[15][15]) );
FA FA_3_143 ( .a(stage_2[15][18]), .b(stage_2[15][19]), .cin(stage_2[15][20]), .cout(stage_3[16][6]), .s(stage_3[15][16]) );
FA FA_3_144 ( .a(stage_2[15][21]), .b(stage_2[15][22]), .cin(stage_2[15][23]), .cout(stage_3[16][7]), .s(stage_3[15][17]) );
FA FA_3_145 ( .a(stage_2[15][24]), .b(stage_2[15][25]), .cin(stage_2[15][26]), .cout(stage_3[16][8]), .s(stage_3[15][18]) );
HA HA_3_12 ( .a(stage_2[15][27]), .b(stage_2[15][28]), .cout(stage_3[16][9]), .s(stage_3[15][19]) );
FA FA_3_146 ( .a(stage_2[16][0]), .b(stage_2[16][1]), .cin(stage_2[16][2]), .cout(stage_3[17][0]), .s(stage_3[16][10]) );
FA FA_3_147 ( .a(stage_2[16][3]), .b(stage_2[16][4]), .cin(stage_2[16][5]), .cout(stage_3[17][1]), .s(stage_3[16][11]) );
FA FA_3_148 ( .a(stage_2[16][6]), .b(stage_2[16][7]), .cin(stage_2[16][8]), .cout(stage_3[17][2]), .s(stage_3[16][12]) );
FA FA_3_149 ( .a(stage_2[16][9]), .b(stage_2[16][10]), .cin(stage_2[16][11]), .cout(stage_3[17][3]), .s(stage_3[16][13]) );
FA FA_3_150 ( .a(stage_2[16][12]), .b(stage_2[16][13]), .cin(stage_2[16][14]), .cout(stage_3[17][4]), .s(stage_3[16][14]) );
FA FA_3_151 ( .a(stage_2[16][15]), .b(stage_2[16][16]), .cin(stage_2[16][17]), .cout(stage_3[17][5]), .s(stage_3[16][15]) );
FA FA_3_152 ( .a(stage_2[16][18]), .b(stage_2[16][19]), .cin(stage_2[16][20]), .cout(stage_3[17][6]), .s(stage_3[16][16]) );
FA FA_3_153 ( .a(stage_2[17][0]), .b(stage_2[17][1]), .cin(stage_2[17][2]), .cout(stage_3[18][0]), .s(stage_3[17][7]) );
FA FA_3_154 ( .a(stage_2[17][3]), .b(stage_2[17][4]), .cin(stage_2[17][5]), .cout(stage_3[18][1]), .s(stage_3[17][8]) );
assign stage_3[17][9] = stage_2[17][6];

wire stage_4 [`NBIT+4:0][`NDATA*2:0];
FA FA_4_0 ( .a(stage_3[0][0]), .b(stage_3[0][1]), .cin(stage_3[0][2]), .cout(stage_4[1][0]), .s(stage_4[0][0]) );
HA HA_4_0 ( .a(stage_3[0][3]), .b(stage_3[0][4]), .cout(stage_4[1][1]), .s(stage_4[0][1]) );
FA FA_4_1 ( .a(stage_3[1][0]), .b(stage_3[1][1]), .cin(stage_3[1][2]), .cout(stage_4[2][0]), .s(stage_4[1][2]) );
FA FA_4_2 ( .a(stage_3[1][3]), .b(stage_3[1][4]), .cin(stage_3[1][5]), .cout(stage_4[2][1]), .s(stage_4[1][3]) );
FA FA_4_3 ( .a(stage_3[1][6]), .b(stage_3[1][7]), .cin(stage_3[1][8]), .cout(stage_4[2][2]), .s(stage_4[1][4]) );
FA FA_4_4 ( .a(stage_3[1][9]), .b(stage_3[1][10]), .cin(stage_3[1][11]), .cout(stage_4[2][3]), .s(stage_4[1][5]) );
FA FA_4_5 ( .a(stage_3[1][12]), .b(stage_3[1][13]), .cin(stage_3[1][14]), .cout(stage_4[2][4]), .s(stage_4[1][6]) );
HA HA_4_1 ( .a(stage_3[1][15]), .b(stage_3[1][16]), .cout(stage_4[2][5]), .s(stage_4[1][7]) );
FA FA_4_6 ( .a(stage_3[2][0]), .b(stage_3[2][1]), .cin(stage_3[2][2]), .cout(stage_4[3][0]), .s(stage_4[2][6]) );
FA FA_4_7 ( .a(stage_3[2][3]), .b(stage_3[2][4]), .cin(stage_3[2][5]), .cout(stage_4[3][1]), .s(stage_4[2][7]) );
FA FA_4_8 ( .a(stage_3[2][6]), .b(stage_3[2][7]), .cin(stage_3[2][8]), .cout(stage_4[3][2]), .s(stage_4[2][8]) );
FA FA_4_9 ( .a(stage_3[2][9]), .b(stage_3[2][10]), .cin(stage_3[2][11]), .cout(stage_4[3][3]), .s(stage_4[2][9]) );
FA FA_4_10 ( .a(stage_3[2][12]), .b(stage_3[2][13]), .cin(stage_3[2][14]), .cout(stage_4[3][4]), .s(stage_4[2][10]) );
FA FA_4_11 ( .a(stage_3[2][15]), .b(stage_3[2][16]), .cin(stage_3[2][17]), .cout(stage_4[3][5]), .s(stage_4[2][11]) );
FA FA_4_12 ( .a(stage_3[2][18]), .b(stage_3[2][19]), .cin(stage_3[2][20]), .cout(stage_4[3][6]), .s(stage_4[2][12]) );
FA FA_4_13 ( .a(stage_3[2][21]), .b(stage_3[2][22]), .cin(stage_3[2][23]), .cout(stage_4[3][7]), .s(stage_4[2][13]) );
assign stage_4[2][14] = stage_3[2][24];
FA FA_4_14 ( .a(stage_3[3][0]), .b(stage_3[3][1]), .cin(stage_3[3][2]), .cout(stage_4[4][0]), .s(stage_4[3][8]) );
FA FA_4_15 ( .a(stage_3[3][3]), .b(stage_3[3][4]), .cin(stage_3[3][5]), .cout(stage_4[4][1]), .s(stage_4[3][9]) );
FA FA_4_16 ( .a(stage_3[3][6]), .b(stage_3[3][7]), .cin(stage_3[3][8]), .cout(stage_4[4][2]), .s(stage_4[3][10]) );
FA FA_4_17 ( .a(stage_3[3][9]), .b(stage_3[3][10]), .cin(stage_3[3][11]), .cout(stage_4[4][3]), .s(stage_4[3][11]) );
FA FA_4_18 ( .a(stage_3[3][12]), .b(stage_3[3][13]), .cin(stage_3[3][14]), .cout(stage_4[4][4]), .s(stage_4[3][12]) );
FA FA_4_19 ( .a(stage_3[3][15]), .b(stage_3[3][16]), .cin(stage_3[3][17]), .cout(stage_4[4][5]), .s(stage_4[3][13]) );
FA FA_4_20 ( .a(stage_3[3][18]), .b(stage_3[3][19]), .cin(stage_3[3][20]), .cout(stage_4[4][6]), .s(stage_4[3][14]) );
assign stage_4[3][15] = stage_3[3][21];
FA FA_4_21 ( .a(stage_3[4][0]), .b(stage_3[4][1]), .cin(stage_3[4][2]), .cout(stage_4[5][0]), .s(stage_4[4][7]) );
FA FA_4_22 ( .a(stage_3[4][3]), .b(stage_3[4][4]), .cin(stage_3[4][5]), .cout(stage_4[5][1]), .s(stage_4[4][8]) );
FA FA_4_23 ( .a(stage_3[4][6]), .b(stage_3[4][7]), .cin(stage_3[4][8]), .cout(stage_4[5][2]), .s(stage_4[4][9]) );
FA FA_4_24 ( .a(stage_3[4][9]), .b(stage_3[4][10]), .cin(stage_3[4][11]), .cout(stage_4[5][3]), .s(stage_4[4][10]) );
FA FA_4_25 ( .a(stage_3[4][12]), .b(stage_3[4][13]), .cin(stage_3[4][14]), .cout(stage_4[5][4]), .s(stage_4[4][11]) );
FA FA_4_26 ( .a(stage_3[4][15]), .b(stage_3[4][16]), .cin(stage_3[4][17]), .cout(stage_4[5][5]), .s(stage_4[4][12]) );
HA HA_4_2 ( .a(stage_3[4][18]), .b(stage_3[4][19]), .cout(stage_4[5][6]), .s(stage_4[4][13]) );
FA FA_4_27 ( .a(stage_3[5][0]), .b(stage_3[5][1]), .cin(stage_3[5][2]), .cout(stage_4[6][0]), .s(stage_4[5][7]) );
FA FA_4_28 ( .a(stage_3[5][3]), .b(stage_3[5][4]), .cin(stage_3[5][5]), .cout(stage_4[6][1]), .s(stage_4[5][8]) );
FA FA_4_29 ( .a(stage_3[5][6]), .b(stage_3[5][7]), .cin(stage_3[5][8]), .cout(stage_4[6][2]), .s(stage_4[5][9]) );
FA FA_4_30 ( .a(stage_3[5][9]), .b(stage_3[5][10]), .cin(stage_3[5][11]), .cout(stage_4[6][3]), .s(stage_4[5][10]) );
FA FA_4_31 ( .a(stage_3[5][12]), .b(stage_3[5][13]), .cin(stage_3[5][14]), .cout(stage_4[6][4]), .s(stage_4[5][11]) );
FA FA_4_32 ( .a(stage_3[5][15]), .b(stage_3[5][16]), .cin(stage_3[5][17]), .cout(stage_4[6][5]), .s(stage_4[5][12]) );
HA HA_4_3 ( .a(stage_3[5][18]), .b(stage_3[5][19]), .cout(stage_4[6][6]), .s(stage_4[5][13]) );
FA FA_4_33 ( .a(stage_3[6][0]), .b(stage_3[6][1]), .cin(stage_3[6][2]), .cout(stage_4[7][0]), .s(stage_4[6][7]) );
FA FA_4_34 ( .a(stage_3[6][3]), .b(stage_3[6][4]), .cin(stage_3[6][5]), .cout(stage_4[7][1]), .s(stage_4[6][8]) );
FA FA_4_35 ( .a(stage_3[6][6]), .b(stage_3[6][7]), .cin(stage_3[6][8]), .cout(stage_4[7][2]), .s(stage_4[6][9]) );
FA FA_4_36 ( .a(stage_3[6][9]), .b(stage_3[6][10]), .cin(stage_3[6][11]), .cout(stage_4[7][3]), .s(stage_4[6][10]) );
FA FA_4_37 ( .a(stage_3[6][12]), .b(stage_3[6][13]), .cin(stage_3[6][14]), .cout(stage_4[7][4]), .s(stage_4[6][11]) );
FA FA_4_38 ( .a(stage_3[6][15]), .b(stage_3[6][16]), .cin(stage_3[6][17]), .cout(stage_4[7][5]), .s(stage_4[6][12]) );
HA HA_4_4 ( .a(stage_3[6][18]), .b(stage_3[6][19]), .cout(stage_4[7][6]), .s(stage_4[6][13]) );
FA FA_4_39 ( .a(stage_3[7][0]), .b(stage_3[7][1]), .cin(stage_3[7][2]), .cout(stage_4[8][0]), .s(stage_4[7][7]) );
FA FA_4_40 ( .a(stage_3[7][3]), .b(stage_3[7][4]), .cin(stage_3[7][5]), .cout(stage_4[8][1]), .s(stage_4[7][8]) );
FA FA_4_41 ( .a(stage_3[7][6]), .b(stage_3[7][7]), .cin(stage_3[7][8]), .cout(stage_4[8][2]), .s(stage_4[7][9]) );
FA FA_4_42 ( .a(stage_3[7][9]), .b(stage_3[7][10]), .cin(stage_3[7][11]), .cout(stage_4[8][3]), .s(stage_4[7][10]) );
FA FA_4_43 ( .a(stage_3[7][12]), .b(stage_3[7][13]), .cin(stage_3[7][14]), .cout(stage_4[8][4]), .s(stage_4[7][11]) );
FA FA_4_44 ( .a(stage_3[7][15]), .b(stage_3[7][16]), .cin(stage_3[7][17]), .cout(stage_4[8][5]), .s(stage_4[7][12]) );
HA HA_4_5 ( .a(stage_3[7][18]), .b(stage_3[7][19]), .cout(stage_4[8][6]), .s(stage_4[7][13]) );
FA FA_4_45 ( .a(stage_3[8][0]), .b(stage_3[8][1]), .cin(stage_3[8][2]), .cout(stage_4[9][0]), .s(stage_4[8][7]) );
FA FA_4_46 ( .a(stage_3[8][3]), .b(stage_3[8][4]), .cin(stage_3[8][5]), .cout(stage_4[9][1]), .s(stage_4[8][8]) );
FA FA_4_47 ( .a(stage_3[8][6]), .b(stage_3[8][7]), .cin(stage_3[8][8]), .cout(stage_4[9][2]), .s(stage_4[8][9]) );
FA FA_4_48 ( .a(stage_3[8][9]), .b(stage_3[8][10]), .cin(stage_3[8][11]), .cout(stage_4[9][3]), .s(stage_4[8][10]) );
FA FA_4_49 ( .a(stage_3[8][12]), .b(stage_3[8][13]), .cin(stage_3[8][14]), .cout(stage_4[9][4]), .s(stage_4[8][11]) );
FA FA_4_50 ( .a(stage_3[8][15]), .b(stage_3[8][16]), .cin(stage_3[8][17]), .cout(stage_4[9][5]), .s(stage_4[8][12]) );
HA HA_4_6 ( .a(stage_3[8][18]), .b(stage_3[8][19]), .cout(stage_4[9][6]), .s(stage_4[8][13]) );
FA FA_4_51 ( .a(stage_3[9][0]), .b(stage_3[9][1]), .cin(stage_3[9][2]), .cout(stage_4[10][0]), .s(stage_4[9][7]) );
FA FA_4_52 ( .a(stage_3[9][3]), .b(stage_3[9][4]), .cin(stage_3[9][5]), .cout(stage_4[10][1]), .s(stage_4[9][8]) );
FA FA_4_53 ( .a(stage_3[9][6]), .b(stage_3[9][7]), .cin(stage_3[9][8]), .cout(stage_4[10][2]), .s(stage_4[9][9]) );
FA FA_4_54 ( .a(stage_3[9][9]), .b(stage_3[9][10]), .cin(stage_3[9][11]), .cout(stage_4[10][3]), .s(stage_4[9][10]) );
FA FA_4_55 ( .a(stage_3[9][12]), .b(stage_3[9][13]), .cin(stage_3[9][14]), .cout(stage_4[10][4]), .s(stage_4[9][11]) );
FA FA_4_56 ( .a(stage_3[9][15]), .b(stage_3[9][16]), .cin(stage_3[9][17]), .cout(stage_4[10][5]), .s(stage_4[9][12]) );
HA HA_4_7 ( .a(stage_3[9][18]), .b(stage_3[9][19]), .cout(stage_4[10][6]), .s(stage_4[9][13]) );
FA FA_4_57 ( .a(stage_3[10][0]), .b(stage_3[10][1]), .cin(stage_3[10][2]), .cout(stage_4[11][0]), .s(stage_4[10][7]) );
FA FA_4_58 ( .a(stage_3[10][3]), .b(stage_3[10][4]), .cin(stage_3[10][5]), .cout(stage_4[11][1]), .s(stage_4[10][8]) );
FA FA_4_59 ( .a(stage_3[10][6]), .b(stage_3[10][7]), .cin(stage_3[10][8]), .cout(stage_4[11][2]), .s(stage_4[10][9]) );
FA FA_4_60 ( .a(stage_3[10][9]), .b(stage_3[10][10]), .cin(stage_3[10][11]), .cout(stage_4[11][3]), .s(stage_4[10][10]) );
FA FA_4_61 ( .a(stage_3[10][12]), .b(stage_3[10][13]), .cin(stage_3[10][14]), .cout(stage_4[11][4]), .s(stage_4[10][11]) );
FA FA_4_62 ( .a(stage_3[10][15]), .b(stage_3[10][16]), .cin(stage_3[10][17]), .cout(stage_4[11][5]), .s(stage_4[10][12]) );
HA HA_4_8 ( .a(stage_3[10][18]), .b(stage_3[10][19]), .cout(stage_4[11][6]), .s(stage_4[10][13]) );
FA FA_4_63 ( .a(stage_3[11][0]), .b(stage_3[11][1]), .cin(stage_3[11][2]), .cout(stage_4[12][0]), .s(stage_4[11][7]) );
FA FA_4_64 ( .a(stage_3[11][3]), .b(stage_3[11][4]), .cin(stage_3[11][5]), .cout(stage_4[12][1]), .s(stage_4[11][8]) );
FA FA_4_65 ( .a(stage_3[11][6]), .b(stage_3[11][7]), .cin(stage_3[11][8]), .cout(stage_4[12][2]), .s(stage_4[11][9]) );
FA FA_4_66 ( .a(stage_3[11][9]), .b(stage_3[11][10]), .cin(stage_3[11][11]), .cout(stage_4[12][3]), .s(stage_4[11][10]) );
FA FA_4_67 ( .a(stage_3[11][12]), .b(stage_3[11][13]), .cin(stage_3[11][14]), .cout(stage_4[12][4]), .s(stage_4[11][11]) );
FA FA_4_68 ( .a(stage_3[11][15]), .b(stage_3[11][16]), .cin(stage_3[11][17]), .cout(stage_4[12][5]), .s(stage_4[11][12]) );
HA HA_4_9 ( .a(stage_3[11][18]), .b(stage_3[11][19]), .cout(stage_4[12][6]), .s(stage_4[11][13]) );
FA FA_4_69 ( .a(stage_3[12][0]), .b(stage_3[12][1]), .cin(stage_3[12][2]), .cout(stage_4[13][0]), .s(stage_4[12][7]) );
FA FA_4_70 ( .a(stage_3[12][3]), .b(stage_3[12][4]), .cin(stage_3[12][5]), .cout(stage_4[13][1]), .s(stage_4[12][8]) );
FA FA_4_71 ( .a(stage_3[12][6]), .b(stage_3[12][7]), .cin(stage_3[12][8]), .cout(stage_4[13][2]), .s(stage_4[12][9]) );
FA FA_4_72 ( .a(stage_3[12][9]), .b(stage_3[12][10]), .cin(stage_3[12][11]), .cout(stage_4[13][3]), .s(stage_4[12][10]) );
FA FA_4_73 ( .a(stage_3[12][12]), .b(stage_3[12][13]), .cin(stage_3[12][14]), .cout(stage_4[13][4]), .s(stage_4[12][11]) );
FA FA_4_74 ( .a(stage_3[12][15]), .b(stage_3[12][16]), .cin(stage_3[12][17]), .cout(stage_4[13][5]), .s(stage_4[12][12]) );
HA HA_4_10 ( .a(stage_3[12][18]), .b(stage_3[12][19]), .cout(stage_4[13][6]), .s(stage_4[12][13]) );
FA FA_4_75 ( .a(stage_3[13][0]), .b(stage_3[13][1]), .cin(stage_3[13][2]), .cout(stage_4[14][0]), .s(stage_4[13][7]) );
FA FA_4_76 ( .a(stage_3[13][3]), .b(stage_3[13][4]), .cin(stage_3[13][5]), .cout(stage_4[14][1]), .s(stage_4[13][8]) );
FA FA_4_77 ( .a(stage_3[13][6]), .b(stage_3[13][7]), .cin(stage_3[13][8]), .cout(stage_4[14][2]), .s(stage_4[13][9]) );
FA FA_4_78 ( .a(stage_3[13][9]), .b(stage_3[13][10]), .cin(stage_3[13][11]), .cout(stage_4[14][3]), .s(stage_4[13][10]) );
FA FA_4_79 ( .a(stage_3[13][12]), .b(stage_3[13][13]), .cin(stage_3[13][14]), .cout(stage_4[14][4]), .s(stage_4[13][11]) );
FA FA_4_80 ( .a(stage_3[13][15]), .b(stage_3[13][16]), .cin(stage_3[13][17]), .cout(stage_4[14][5]), .s(stage_4[13][12]) );
HA HA_4_11 ( .a(stage_3[13][18]), .b(stage_3[13][19]), .cout(stage_4[14][6]), .s(stage_4[13][13]) );
FA FA_4_81 ( .a(stage_3[14][0]), .b(stage_3[14][1]), .cin(stage_3[14][2]), .cout(stage_4[15][0]), .s(stage_4[14][7]) );
FA FA_4_82 ( .a(stage_3[14][3]), .b(stage_3[14][4]), .cin(stage_3[14][5]), .cout(stage_4[15][1]), .s(stage_4[14][8]) );
FA FA_4_83 ( .a(stage_3[14][6]), .b(stage_3[14][7]), .cin(stage_3[14][8]), .cout(stage_4[15][2]), .s(stage_4[14][9]) );
FA FA_4_84 ( .a(stage_3[14][9]), .b(stage_3[14][10]), .cin(stage_3[14][11]), .cout(stage_4[15][3]), .s(stage_4[14][10]) );
FA FA_4_85 ( .a(stage_3[14][12]), .b(stage_3[14][13]), .cin(stage_3[14][14]), .cout(stage_4[15][4]), .s(stage_4[14][11]) );
FA FA_4_86 ( .a(stage_3[14][15]), .b(stage_3[14][16]), .cin(stage_3[14][17]), .cout(stage_4[15][5]), .s(stage_4[14][12]) );
HA HA_4_12 ( .a(stage_3[14][18]), .b(stage_3[14][19]), .cout(stage_4[15][6]), .s(stage_4[14][13]) );
FA FA_4_87 ( .a(stage_3[15][0]), .b(stage_3[15][1]), .cin(stage_3[15][2]), .cout(stage_4[16][0]), .s(stage_4[15][7]) );
FA FA_4_88 ( .a(stage_3[15][3]), .b(stage_3[15][4]), .cin(stage_3[15][5]), .cout(stage_4[16][1]), .s(stage_4[15][8]) );
FA FA_4_89 ( .a(stage_3[15][6]), .b(stage_3[15][7]), .cin(stage_3[15][8]), .cout(stage_4[16][2]), .s(stage_4[15][9]) );
FA FA_4_90 ( .a(stage_3[15][9]), .b(stage_3[15][10]), .cin(stage_3[15][11]), .cout(stage_4[16][3]), .s(stage_4[15][10]) );
FA FA_4_91 ( .a(stage_3[15][12]), .b(stage_3[15][13]), .cin(stage_3[15][14]), .cout(stage_4[16][4]), .s(stage_4[15][11]) );
FA FA_4_92 ( .a(stage_3[15][15]), .b(stage_3[15][16]), .cin(stage_3[15][17]), .cout(stage_4[16][5]), .s(stage_4[15][12]) );
HA HA_4_13 ( .a(stage_3[15][18]), .b(stage_3[15][19]), .cout(stage_4[16][6]), .s(stage_4[15][13]) );
FA FA_4_93 ( .a(stage_3[16][0]), .b(stage_3[16][1]), .cin(stage_3[16][2]), .cout(stage_4[17][0]), .s(stage_4[16][7]) );
FA FA_4_94 ( .a(stage_3[16][3]), .b(stage_3[16][4]), .cin(stage_3[16][5]), .cout(stage_4[17][1]), .s(stage_4[16][8]) );
FA FA_4_95 ( .a(stage_3[16][6]), .b(stage_3[16][7]), .cin(stage_3[16][8]), .cout(stage_4[17][2]), .s(stage_4[16][9]) );
FA FA_4_96 ( .a(stage_3[16][9]), .b(stage_3[16][10]), .cin(stage_3[16][11]), .cout(stage_4[17][3]), .s(stage_4[16][10]) );
FA FA_4_97 ( .a(stage_3[16][12]), .b(stage_3[16][13]), .cin(stage_3[16][14]), .cout(stage_4[17][4]), .s(stage_4[16][11]) );
HA HA_4_14 ( .a(stage_3[16][15]), .b(stage_3[16][16]), .cout(stage_4[17][5]), .s(stage_4[16][12]) );
FA FA_4_98 ( .a(stage_3[17][0]), .b(stage_3[17][1]), .cin(stage_3[17][2]), .cout(stage_4[18][0]), .s(stage_4[17][6]) );
FA FA_4_99 ( .a(stage_3[17][3]), .b(stage_3[17][4]), .cin(stage_3[17][5]), .cout(stage_4[18][1]), .s(stage_4[17][7]) );
FA FA_4_100 ( .a(stage_3[17][6]), .b(stage_3[17][7]), .cin(stage_3[17][8]), .cout(stage_4[18][2]), .s(stage_4[17][8]) );
assign stage_4[17][9] = stage_3[17][9];
HA HA_4_15 ( .a(stage_3[18][0]), .b(stage_3[18][1]), .cout(stage_4[19][0]), .s(stage_4[18][3]) );

wire stage_5 [`NBIT+5:0][`NDATA*2:0];
HA HA_5_0 ( .a(stage_4[0][0]), .b(stage_4[0][1]), .cout(stage_5[1][0]), .s(stage_5[0][0]) );
FA FA_5_0 ( .a(stage_4[1][0]), .b(stage_4[1][1]), .cin(stage_4[1][2]), .cout(stage_5[2][0]), .s(stage_5[1][1]) );
FA FA_5_1 ( .a(stage_4[1][3]), .b(stage_4[1][4]), .cin(stage_4[1][5]), .cout(stage_5[2][1]), .s(stage_5[1][2]) );
HA HA_5_1 ( .a(stage_4[1][6]), .b(stage_4[1][7]), .cout(stage_5[2][2]), .s(stage_5[1][3]) );
FA FA_5_2 ( .a(stage_4[2][0]), .b(stage_4[2][1]), .cin(stage_4[2][2]), .cout(stage_5[3][0]), .s(stage_5[2][3]) );
FA FA_5_3 ( .a(stage_4[2][3]), .b(stage_4[2][4]), .cin(stage_4[2][5]), .cout(stage_5[3][1]), .s(stage_5[2][4]) );
FA FA_5_4 ( .a(stage_4[2][6]), .b(stage_4[2][7]), .cin(stage_4[2][8]), .cout(stage_5[3][2]), .s(stage_5[2][5]) );
FA FA_5_5 ( .a(stage_4[2][9]), .b(stage_4[2][10]), .cin(stage_4[2][11]), .cout(stage_5[3][3]), .s(stage_5[2][6]) );
FA FA_5_6 ( .a(stage_4[2][12]), .b(stage_4[2][13]), .cin(stage_4[2][14]), .cout(stage_5[3][4]), .s(stage_5[2][7]) );
FA FA_5_7 ( .a(stage_4[3][0]), .b(stage_4[3][1]), .cin(stage_4[3][2]), .cout(stage_5[4][0]), .s(stage_5[3][5]) );
FA FA_5_8 ( .a(stage_4[3][3]), .b(stage_4[3][4]), .cin(stage_4[3][5]), .cout(stage_5[4][1]), .s(stage_5[3][6]) );
FA FA_5_9 ( .a(stage_4[3][6]), .b(stage_4[3][7]), .cin(stage_4[3][8]), .cout(stage_5[4][2]), .s(stage_5[3][7]) );
FA FA_5_10 ( .a(stage_4[3][9]), .b(stage_4[3][10]), .cin(stage_4[3][11]), .cout(stage_5[4][3]), .s(stage_5[3][8]) );
FA FA_5_11 ( .a(stage_4[3][12]), .b(stage_4[3][13]), .cin(stage_4[3][14]), .cout(stage_5[4][4]), .s(stage_5[3][9]) );
assign stage_5[3][10] = stage_4[3][15];
FA FA_5_12 ( .a(stage_4[4][0]), .b(stage_4[4][1]), .cin(stage_4[4][2]), .cout(stage_5[5][0]), .s(stage_5[4][5]) );
FA FA_5_13 ( .a(stage_4[4][3]), .b(stage_4[4][4]), .cin(stage_4[4][5]), .cout(stage_5[5][1]), .s(stage_5[4][6]) );
FA FA_5_14 ( .a(stage_4[4][6]), .b(stage_4[4][7]), .cin(stage_4[4][8]), .cout(stage_5[5][2]), .s(stage_5[4][7]) );
FA FA_5_15 ( .a(stage_4[4][9]), .b(stage_4[4][10]), .cin(stage_4[4][11]), .cout(stage_5[5][3]), .s(stage_5[4][8]) );
HA HA_5_2 ( .a(stage_4[4][12]), .b(stage_4[4][13]), .cout(stage_5[5][4]), .s(stage_5[4][9]) );
FA FA_5_16 ( .a(stage_4[5][0]), .b(stage_4[5][1]), .cin(stage_4[5][2]), .cout(stage_5[6][0]), .s(stage_5[5][5]) );
FA FA_5_17 ( .a(stage_4[5][3]), .b(stage_4[5][4]), .cin(stage_4[5][5]), .cout(stage_5[6][1]), .s(stage_5[5][6]) );
FA FA_5_18 ( .a(stage_4[5][6]), .b(stage_4[5][7]), .cin(stage_4[5][8]), .cout(stage_5[6][2]), .s(stage_5[5][7]) );
FA FA_5_19 ( .a(stage_4[5][9]), .b(stage_4[5][10]), .cin(stage_4[5][11]), .cout(stage_5[6][3]), .s(stage_5[5][8]) );
HA HA_5_3 ( .a(stage_4[5][12]), .b(stage_4[5][13]), .cout(stage_5[6][4]), .s(stage_5[5][9]) );
FA FA_5_20 ( .a(stage_4[6][0]), .b(stage_4[6][1]), .cin(stage_4[6][2]), .cout(stage_5[7][0]), .s(stage_5[6][5]) );
FA FA_5_21 ( .a(stage_4[6][3]), .b(stage_4[6][4]), .cin(stage_4[6][5]), .cout(stage_5[7][1]), .s(stage_5[6][6]) );
FA FA_5_22 ( .a(stage_4[6][6]), .b(stage_4[6][7]), .cin(stage_4[6][8]), .cout(stage_5[7][2]), .s(stage_5[6][7]) );
FA FA_5_23 ( .a(stage_4[6][9]), .b(stage_4[6][10]), .cin(stage_4[6][11]), .cout(stage_5[7][3]), .s(stage_5[6][8]) );
HA HA_5_4 ( .a(stage_4[6][12]), .b(stage_4[6][13]), .cout(stage_5[7][4]), .s(stage_5[6][9]) );
FA FA_5_24 ( .a(stage_4[7][0]), .b(stage_4[7][1]), .cin(stage_4[7][2]), .cout(stage_5[8][0]), .s(stage_5[7][5]) );
FA FA_5_25 ( .a(stage_4[7][3]), .b(stage_4[7][4]), .cin(stage_4[7][5]), .cout(stage_5[8][1]), .s(stage_5[7][6]) );
FA FA_5_26 ( .a(stage_4[7][6]), .b(stage_4[7][7]), .cin(stage_4[7][8]), .cout(stage_5[8][2]), .s(stage_5[7][7]) );
FA FA_5_27 ( .a(stage_4[7][9]), .b(stage_4[7][10]), .cin(stage_4[7][11]), .cout(stage_5[8][3]), .s(stage_5[7][8]) );
HA HA_5_5 ( .a(stage_4[7][12]), .b(stage_4[7][13]), .cout(stage_5[8][4]), .s(stage_5[7][9]) );
FA FA_5_28 ( .a(stage_4[8][0]), .b(stage_4[8][1]), .cin(stage_4[8][2]), .cout(stage_5[9][0]), .s(stage_5[8][5]) );
FA FA_5_29 ( .a(stage_4[8][3]), .b(stage_4[8][4]), .cin(stage_4[8][5]), .cout(stage_5[9][1]), .s(stage_5[8][6]) );
FA FA_5_30 ( .a(stage_4[8][6]), .b(stage_4[8][7]), .cin(stage_4[8][8]), .cout(stage_5[9][2]), .s(stage_5[8][7]) );
FA FA_5_31 ( .a(stage_4[8][9]), .b(stage_4[8][10]), .cin(stage_4[8][11]), .cout(stage_5[9][3]), .s(stage_5[8][8]) );
HA HA_5_6 ( .a(stage_4[8][12]), .b(stage_4[8][13]), .cout(stage_5[9][4]), .s(stage_5[8][9]) );
FA FA_5_32 ( .a(stage_4[9][0]), .b(stage_4[9][1]), .cin(stage_4[9][2]), .cout(stage_5[10][0]), .s(stage_5[9][5]) );
FA FA_5_33 ( .a(stage_4[9][3]), .b(stage_4[9][4]), .cin(stage_4[9][5]), .cout(stage_5[10][1]), .s(stage_5[9][6]) );
FA FA_5_34 ( .a(stage_4[9][6]), .b(stage_4[9][7]), .cin(stage_4[9][8]), .cout(stage_5[10][2]), .s(stage_5[9][7]) );
FA FA_5_35 ( .a(stage_4[9][9]), .b(stage_4[9][10]), .cin(stage_4[9][11]), .cout(stage_5[10][3]), .s(stage_5[9][8]) );
HA HA_5_7 ( .a(stage_4[9][12]), .b(stage_4[9][13]), .cout(stage_5[10][4]), .s(stage_5[9][9]) );
FA FA_5_36 ( .a(stage_4[10][0]), .b(stage_4[10][1]), .cin(stage_4[10][2]), .cout(stage_5[11][0]), .s(stage_5[10][5]) );
FA FA_5_37 ( .a(stage_4[10][3]), .b(stage_4[10][4]), .cin(stage_4[10][5]), .cout(stage_5[11][1]), .s(stage_5[10][6]) );
FA FA_5_38 ( .a(stage_4[10][6]), .b(stage_4[10][7]), .cin(stage_4[10][8]), .cout(stage_5[11][2]), .s(stage_5[10][7]) );
FA FA_5_39 ( .a(stage_4[10][9]), .b(stage_4[10][10]), .cin(stage_4[10][11]), .cout(stage_5[11][3]), .s(stage_5[10][8]) );
HA HA_5_8 ( .a(stage_4[10][12]), .b(stage_4[10][13]), .cout(stage_5[11][4]), .s(stage_5[10][9]) );
FA FA_5_40 ( .a(stage_4[11][0]), .b(stage_4[11][1]), .cin(stage_4[11][2]), .cout(stage_5[12][0]), .s(stage_5[11][5]) );
FA FA_5_41 ( .a(stage_4[11][3]), .b(stage_4[11][4]), .cin(stage_4[11][5]), .cout(stage_5[12][1]), .s(stage_5[11][6]) );
FA FA_5_42 ( .a(stage_4[11][6]), .b(stage_4[11][7]), .cin(stage_4[11][8]), .cout(stage_5[12][2]), .s(stage_5[11][7]) );
FA FA_5_43 ( .a(stage_4[11][9]), .b(stage_4[11][10]), .cin(stage_4[11][11]), .cout(stage_5[12][3]), .s(stage_5[11][8]) );
HA HA_5_9 ( .a(stage_4[11][12]), .b(stage_4[11][13]), .cout(stage_5[12][4]), .s(stage_5[11][9]) );
FA FA_5_44 ( .a(stage_4[12][0]), .b(stage_4[12][1]), .cin(stage_4[12][2]), .cout(stage_5[13][0]), .s(stage_5[12][5]) );
FA FA_5_45 ( .a(stage_4[12][3]), .b(stage_4[12][4]), .cin(stage_4[12][5]), .cout(stage_5[13][1]), .s(stage_5[12][6]) );
FA FA_5_46 ( .a(stage_4[12][6]), .b(stage_4[12][7]), .cin(stage_4[12][8]), .cout(stage_5[13][2]), .s(stage_5[12][7]) );
FA FA_5_47 ( .a(stage_4[12][9]), .b(stage_4[12][10]), .cin(stage_4[12][11]), .cout(stage_5[13][3]), .s(stage_5[12][8]) );
HA HA_5_10 ( .a(stage_4[12][12]), .b(stage_4[12][13]), .cout(stage_5[13][4]), .s(stage_5[12][9]) );
FA FA_5_48 ( .a(stage_4[13][0]), .b(stage_4[13][1]), .cin(stage_4[13][2]), .cout(stage_5[14][0]), .s(stage_5[13][5]) );
FA FA_5_49 ( .a(stage_4[13][3]), .b(stage_4[13][4]), .cin(stage_4[13][5]), .cout(stage_5[14][1]), .s(stage_5[13][6]) );
FA FA_5_50 ( .a(stage_4[13][6]), .b(stage_4[13][7]), .cin(stage_4[13][8]), .cout(stage_5[14][2]), .s(stage_5[13][7]) );
FA FA_5_51 ( .a(stage_4[13][9]), .b(stage_4[13][10]), .cin(stage_4[13][11]), .cout(stage_5[14][3]), .s(stage_5[13][8]) );
HA HA_5_11 ( .a(stage_4[13][12]), .b(stage_4[13][13]), .cout(stage_5[14][4]), .s(stage_5[13][9]) );
FA FA_5_52 ( .a(stage_4[14][0]), .b(stage_4[14][1]), .cin(stage_4[14][2]), .cout(stage_5[15][0]), .s(stage_5[14][5]) );
FA FA_5_53 ( .a(stage_4[14][3]), .b(stage_4[14][4]), .cin(stage_4[14][5]), .cout(stage_5[15][1]), .s(stage_5[14][6]) );
FA FA_5_54 ( .a(stage_4[14][6]), .b(stage_4[14][7]), .cin(stage_4[14][8]), .cout(stage_5[15][2]), .s(stage_5[14][7]) );
FA FA_5_55 ( .a(stage_4[14][9]), .b(stage_4[14][10]), .cin(stage_4[14][11]), .cout(stage_5[15][3]), .s(stage_5[14][8]) );
HA HA_5_12 ( .a(stage_4[14][12]), .b(stage_4[14][13]), .cout(stage_5[15][4]), .s(stage_5[14][9]) );
FA FA_5_56 ( .a(stage_4[15][0]), .b(stage_4[15][1]), .cin(stage_4[15][2]), .cout(stage_5[16][0]), .s(stage_5[15][5]) );
FA FA_5_57 ( .a(stage_4[15][3]), .b(stage_4[15][4]), .cin(stage_4[15][5]), .cout(stage_5[16][1]), .s(stage_5[15][6]) );
FA FA_5_58 ( .a(stage_4[15][6]), .b(stage_4[15][7]), .cin(stage_4[15][8]), .cout(stage_5[16][2]), .s(stage_5[15][7]) );
FA FA_5_59 ( .a(stage_4[15][9]), .b(stage_4[15][10]), .cin(stage_4[15][11]), .cout(stage_5[16][3]), .s(stage_5[15][8]) );
HA HA_5_13 ( .a(stage_4[15][12]), .b(stage_4[15][13]), .cout(stage_5[16][4]), .s(stage_5[15][9]) );
FA FA_5_60 ( .a(stage_4[16][0]), .b(stage_4[16][1]), .cin(stage_4[16][2]), .cout(stage_5[17][0]), .s(stage_5[16][5]) );
FA FA_5_61 ( .a(stage_4[16][3]), .b(stage_4[16][4]), .cin(stage_4[16][5]), .cout(stage_5[17][1]), .s(stage_5[16][6]) );
FA FA_5_62 ( .a(stage_4[16][6]), .b(stage_4[16][7]), .cin(stage_4[16][8]), .cout(stage_5[17][2]), .s(stage_5[16][7]) );
FA FA_5_63 ( .a(stage_4[16][9]), .b(stage_4[16][10]), .cin(stage_4[16][11]), .cout(stage_5[17][3]), .s(stage_5[16][8]) );
assign stage_5[16][9] = stage_4[16][12];
FA FA_5_64 ( .a(stage_4[17][0]), .b(stage_4[17][1]), .cin(stage_4[17][2]), .cout(stage_5[18][0]), .s(stage_5[17][4]) );
FA FA_5_65 ( .a(stage_4[17][3]), .b(stage_4[17][4]), .cin(stage_4[17][5]), .cout(stage_5[18][1]), .s(stage_5[17][5]) );
FA FA_5_66 ( .a(stage_4[17][6]), .b(stage_4[17][7]), .cin(stage_4[17][8]), .cout(stage_5[18][2]), .s(stage_5[17][6]) );
assign stage_5[17][7] = stage_4[17][9];
FA FA_5_67 ( .a(stage_4[18][0]), .b(stage_4[18][1]), .cin(stage_4[18][2]), .cout(stage_5[19][0]), .s(stage_5[18][3]) );
assign stage_5[18][4] = stage_4[18][3];
assign stage_5[19][1] = stage_4[19][0];

wire stage_6 [`NBIT+6:0][`NDATA*2:0];
assign stage_6[0][0] = stage_5[0][0];
FA FA_6_0 ( .a(stage_5[1][0]), .b(stage_5[1][1]), .cin(stage_5[1][2]), .cout(stage_6[2][0]), .s(stage_6[1][0]) );
assign stage_6[1][1] = stage_5[1][3];
FA FA_6_1 ( .a(stage_5[2][0]), .b(stage_5[2][1]), .cin(stage_5[2][2]), .cout(stage_6[3][0]), .s(stage_6[2][1]) );
FA FA_6_2 ( .a(stage_5[2][3]), .b(stage_5[2][4]), .cin(stage_5[2][5]), .cout(stage_6[3][1]), .s(stage_6[2][2]) );
HA HA_6_0 ( .a(stage_5[2][6]), .b(stage_5[2][7]), .cout(stage_6[3][2]), .s(stage_6[2][3]) );
FA FA_6_3 ( .a(stage_5[3][0]), .b(stage_5[3][1]), .cin(stage_5[3][2]), .cout(stage_6[4][0]), .s(stage_6[3][3]) );
FA FA_6_4 ( .a(stage_5[3][3]), .b(stage_5[3][4]), .cin(stage_5[3][5]), .cout(stage_6[4][1]), .s(stage_6[3][4]) );
FA FA_6_5 ( .a(stage_5[3][6]), .b(stage_5[3][7]), .cin(stage_5[3][8]), .cout(stage_6[4][2]), .s(stage_6[3][5]) );
HA HA_6_1 ( .a(stage_5[3][9]), .b(stage_5[3][10]), .cout(stage_6[4][3]), .s(stage_6[3][6]) );
FA FA_6_6 ( .a(stage_5[4][0]), .b(stage_5[4][1]), .cin(stage_5[4][2]), .cout(stage_6[5][0]), .s(stage_6[4][4]) );
FA FA_6_7 ( .a(stage_5[4][3]), .b(stage_5[4][4]), .cin(stage_5[4][5]), .cout(stage_6[5][1]), .s(stage_6[4][5]) );
FA FA_6_8 ( .a(stage_5[4][6]), .b(stage_5[4][7]), .cin(stage_5[4][8]), .cout(stage_6[5][2]), .s(stage_6[4][6]) );
assign stage_6[4][7] = stage_5[4][9];
FA FA_6_9 ( .a(stage_5[5][0]), .b(stage_5[5][1]), .cin(stage_5[5][2]), .cout(stage_6[6][0]), .s(stage_6[5][3]) );
FA FA_6_10 ( .a(stage_5[5][3]), .b(stage_5[5][4]), .cin(stage_5[5][5]), .cout(stage_6[6][1]), .s(stage_6[5][4]) );
FA FA_6_11 ( .a(stage_5[5][6]), .b(stage_5[5][7]), .cin(stage_5[5][8]), .cout(stage_6[6][2]), .s(stage_6[5][5]) );
assign stage_6[5][6] = stage_5[5][9];
FA FA_6_12 ( .a(stage_5[6][0]), .b(stage_5[6][1]), .cin(stage_5[6][2]), .cout(stage_6[7][0]), .s(stage_6[6][3]) );
FA FA_6_13 ( .a(stage_5[6][3]), .b(stage_5[6][4]), .cin(stage_5[6][5]), .cout(stage_6[7][1]), .s(stage_6[6][4]) );
FA FA_6_14 ( .a(stage_5[6][6]), .b(stage_5[6][7]), .cin(stage_5[6][8]), .cout(stage_6[7][2]), .s(stage_6[6][5]) );
assign stage_6[6][6] = stage_5[6][9];
FA FA_6_15 ( .a(stage_5[7][0]), .b(stage_5[7][1]), .cin(stage_5[7][2]), .cout(stage_6[8][0]), .s(stage_6[7][3]) );
FA FA_6_16 ( .a(stage_5[7][3]), .b(stage_5[7][4]), .cin(stage_5[7][5]), .cout(stage_6[8][1]), .s(stage_6[7][4]) );
FA FA_6_17 ( .a(stage_5[7][6]), .b(stage_5[7][7]), .cin(stage_5[7][8]), .cout(stage_6[8][2]), .s(stage_6[7][5]) );
assign stage_6[7][6] = stage_5[7][9];
FA FA_6_18 ( .a(stage_5[8][0]), .b(stage_5[8][1]), .cin(stage_5[8][2]), .cout(stage_6[9][0]), .s(stage_6[8][3]) );
FA FA_6_19 ( .a(stage_5[8][3]), .b(stage_5[8][4]), .cin(stage_5[8][5]), .cout(stage_6[9][1]), .s(stage_6[8][4]) );
FA FA_6_20 ( .a(stage_5[8][6]), .b(stage_5[8][7]), .cin(stage_5[8][8]), .cout(stage_6[9][2]), .s(stage_6[8][5]) );
assign stage_6[8][6] = stage_5[8][9];
FA FA_6_21 ( .a(stage_5[9][0]), .b(stage_5[9][1]), .cin(stage_5[9][2]), .cout(stage_6[10][0]), .s(stage_6[9][3]) );
FA FA_6_22 ( .a(stage_5[9][3]), .b(stage_5[9][4]), .cin(stage_5[9][5]), .cout(stage_6[10][1]), .s(stage_6[9][4]) );
FA FA_6_23 ( .a(stage_5[9][6]), .b(stage_5[9][7]), .cin(stage_5[9][8]), .cout(stage_6[10][2]), .s(stage_6[9][5]) );
assign stage_6[9][6] = stage_5[9][9];
FA FA_6_24 ( .a(stage_5[10][0]), .b(stage_5[10][1]), .cin(stage_5[10][2]), .cout(stage_6[11][0]), .s(stage_6[10][3]) );
FA FA_6_25 ( .a(stage_5[10][3]), .b(stage_5[10][4]), .cin(stage_5[10][5]), .cout(stage_6[11][1]), .s(stage_6[10][4]) );
FA FA_6_26 ( .a(stage_5[10][6]), .b(stage_5[10][7]), .cin(stage_5[10][8]), .cout(stage_6[11][2]), .s(stage_6[10][5]) );
assign stage_6[10][6] = stage_5[10][9];
FA FA_6_27 ( .a(stage_5[11][0]), .b(stage_5[11][1]), .cin(stage_5[11][2]), .cout(stage_6[12][0]), .s(stage_6[11][3]) );
FA FA_6_28 ( .a(stage_5[11][3]), .b(stage_5[11][4]), .cin(stage_5[11][5]), .cout(stage_6[12][1]), .s(stage_6[11][4]) );
FA FA_6_29 ( .a(stage_5[11][6]), .b(stage_5[11][7]), .cin(stage_5[11][8]), .cout(stage_6[12][2]), .s(stage_6[11][5]) );
assign stage_6[11][6] = stage_5[11][9];
FA FA_6_30 ( .a(stage_5[12][0]), .b(stage_5[12][1]), .cin(stage_5[12][2]), .cout(stage_6[13][0]), .s(stage_6[12][3]) );
FA FA_6_31 ( .a(stage_5[12][3]), .b(stage_5[12][4]), .cin(stage_5[12][5]), .cout(stage_6[13][1]), .s(stage_6[12][4]) );
FA FA_6_32 ( .a(stage_5[12][6]), .b(stage_5[12][7]), .cin(stage_5[12][8]), .cout(stage_6[13][2]), .s(stage_6[12][5]) );
assign stage_6[12][6] = stage_5[12][9];
FA FA_6_33 ( .a(stage_5[13][0]), .b(stage_5[13][1]), .cin(stage_5[13][2]), .cout(stage_6[14][0]), .s(stage_6[13][3]) );
FA FA_6_34 ( .a(stage_5[13][3]), .b(stage_5[13][4]), .cin(stage_5[13][5]), .cout(stage_6[14][1]), .s(stage_6[13][4]) );
FA FA_6_35 ( .a(stage_5[13][6]), .b(stage_5[13][7]), .cin(stage_5[13][8]), .cout(stage_6[14][2]), .s(stage_6[13][5]) );
assign stage_6[13][6] = stage_5[13][9];
FA FA_6_36 ( .a(stage_5[14][0]), .b(stage_5[14][1]), .cin(stage_5[14][2]), .cout(stage_6[15][0]), .s(stage_6[14][3]) );
FA FA_6_37 ( .a(stage_5[14][3]), .b(stage_5[14][4]), .cin(stage_5[14][5]), .cout(stage_6[15][1]), .s(stage_6[14][4]) );
FA FA_6_38 ( .a(stage_5[14][6]), .b(stage_5[14][7]), .cin(stage_5[14][8]), .cout(stage_6[15][2]), .s(stage_6[14][5]) );
assign stage_6[14][6] = stage_5[14][9];
FA FA_6_39 ( .a(stage_5[15][0]), .b(stage_5[15][1]), .cin(stage_5[15][2]), .cout(stage_6[16][0]), .s(stage_6[15][3]) );
FA FA_6_40 ( .a(stage_5[15][3]), .b(stage_5[15][4]), .cin(stage_5[15][5]), .cout(stage_6[16][1]), .s(stage_6[15][4]) );
FA FA_6_41 ( .a(stage_5[15][6]), .b(stage_5[15][7]), .cin(stage_5[15][8]), .cout(stage_6[16][2]), .s(stage_6[15][5]) );
assign stage_6[15][6] = stage_5[15][9];
FA FA_6_42 ( .a(stage_5[16][0]), .b(stage_5[16][1]), .cin(stage_5[16][2]), .cout(stage_6[17][0]), .s(stage_6[16][3]) );
FA FA_6_43 ( .a(stage_5[16][3]), .b(stage_5[16][4]), .cin(stage_5[16][5]), .cout(stage_6[17][1]), .s(stage_6[16][4]) );
FA FA_6_44 ( .a(stage_5[16][6]), .b(stage_5[16][7]), .cin(stage_5[16][8]), .cout(stage_6[17][2]), .s(stage_6[16][5]) );
assign stage_6[16][6] = stage_5[16][9];
FA FA_6_45 ( .a(stage_5[17][0]), .b(stage_5[17][1]), .cin(stage_5[17][2]), .cout(stage_6[18][0]), .s(stage_6[17][3]) );
FA FA_6_46 ( .a(stage_5[17][3]), .b(stage_5[17][4]), .cin(stage_5[17][5]), .cout(stage_6[18][1]), .s(stage_6[17][4]) );
HA HA_6_2 ( .a(stage_5[17][6]), .b(stage_5[17][7]), .cout(stage_6[18][2]), .s(stage_6[17][5]) );
FA FA_6_47 ( .a(stage_5[18][0]), .b(stage_5[18][1]), .cin(stage_5[18][2]), .cout(stage_6[19][0]), .s(stage_6[18][3]) );
HA HA_6_3 ( .a(stage_5[18][3]), .b(stage_5[18][4]), .cout(stage_6[19][1]), .s(stage_6[18][4]) );
HA HA_6_4 ( .a(stage_5[19][0]), .b(stage_5[19][1]), .cout(stage_6[20][0]), .s(stage_6[19][2]) );

wire stage_7 [`NBIT+7:0][`NDATA*2:0];
assign stage_7[0][0] = stage_6[0][0];
HA HA_7_0 ( .a(stage_6[1][0]), .b(stage_6[1][1]), .cout(stage_7[2][0]), .s(stage_7[1][0]) );
FA FA_7_0 ( .a(stage_6[2][0]), .b(stage_6[2][1]), .cin(stage_6[2][2]), .cout(stage_7[3][0]), .s(stage_7[2][1]) );
assign stage_7[2][2] = stage_6[2][3];
FA FA_7_1 ( .a(stage_6[3][0]), .b(stage_6[3][1]), .cin(stage_6[3][2]), .cout(stage_7[4][0]), .s(stage_7[3][1]) );
FA FA_7_2 ( .a(stage_6[3][3]), .b(stage_6[3][4]), .cin(stage_6[3][5]), .cout(stage_7[4][1]), .s(stage_7[3][2]) );
assign stage_7[3][3] = stage_6[3][6];
FA FA_7_3 ( .a(stage_6[4][0]), .b(stage_6[4][1]), .cin(stage_6[4][2]), .cout(stage_7[5][0]), .s(stage_7[4][2]) );
FA FA_7_4 ( .a(stage_6[4][3]), .b(stage_6[4][4]), .cin(stage_6[4][5]), .cout(stage_7[5][1]), .s(stage_7[4][3]) );
HA HA_7_1 ( .a(stage_6[4][6]), .b(stage_6[4][7]), .cout(stage_7[5][2]), .s(stage_7[4][4]) );
FA FA_7_5 ( .a(stage_6[5][0]), .b(stage_6[5][1]), .cin(stage_6[5][2]), .cout(stage_7[6][0]), .s(stage_7[5][3]) );
FA FA_7_6 ( .a(stage_6[5][3]), .b(stage_6[5][4]), .cin(stage_6[5][5]), .cout(stage_7[6][1]), .s(stage_7[5][4]) );
assign stage_7[5][5] = stage_6[5][6];
FA FA_7_7 ( .a(stage_6[6][0]), .b(stage_6[6][1]), .cin(stage_6[6][2]), .cout(stage_7[7][0]), .s(stage_7[6][2]) );
FA FA_7_8 ( .a(stage_6[6][3]), .b(stage_6[6][4]), .cin(stage_6[6][5]), .cout(stage_7[7][1]), .s(stage_7[6][3]) );
assign stage_7[6][4] = stage_6[6][6];
FA FA_7_9 ( .a(stage_6[7][0]), .b(stage_6[7][1]), .cin(stage_6[7][2]), .cout(stage_7[8][0]), .s(stage_7[7][2]) );
FA FA_7_10 ( .a(stage_6[7][3]), .b(stage_6[7][4]), .cin(stage_6[7][5]), .cout(stage_7[8][1]), .s(stage_7[7][3]) );
assign stage_7[7][4] = stage_6[7][6];
FA FA_7_11 ( .a(stage_6[8][0]), .b(stage_6[8][1]), .cin(stage_6[8][2]), .cout(stage_7[9][0]), .s(stage_7[8][2]) );
FA FA_7_12 ( .a(stage_6[8][3]), .b(stage_6[8][4]), .cin(stage_6[8][5]), .cout(stage_7[9][1]), .s(stage_7[8][3]) );
assign stage_7[8][4] = stage_6[8][6];
FA FA_7_13 ( .a(stage_6[9][0]), .b(stage_6[9][1]), .cin(stage_6[9][2]), .cout(stage_7[10][0]), .s(stage_7[9][2]) );
FA FA_7_14 ( .a(stage_6[9][3]), .b(stage_6[9][4]), .cin(stage_6[9][5]), .cout(stage_7[10][1]), .s(stage_7[9][3]) );
assign stage_7[9][4] = stage_6[9][6];
FA FA_7_15 ( .a(stage_6[10][0]), .b(stage_6[10][1]), .cin(stage_6[10][2]), .cout(stage_7[11][0]), .s(stage_7[10][2]) );
FA FA_7_16 ( .a(stage_6[10][3]), .b(stage_6[10][4]), .cin(stage_6[10][5]), .cout(stage_7[11][1]), .s(stage_7[10][3]) );
assign stage_7[10][4] = stage_6[10][6];
FA FA_7_17 ( .a(stage_6[11][0]), .b(stage_6[11][1]), .cin(stage_6[11][2]), .cout(stage_7[12][0]), .s(stage_7[11][2]) );
FA FA_7_18 ( .a(stage_6[11][3]), .b(stage_6[11][4]), .cin(stage_6[11][5]), .cout(stage_7[12][1]), .s(stage_7[11][3]) );
assign stage_7[11][4] = stage_6[11][6];
FA FA_7_19 ( .a(stage_6[12][0]), .b(stage_6[12][1]), .cin(stage_6[12][2]), .cout(stage_7[13][0]), .s(stage_7[12][2]) );
FA FA_7_20 ( .a(stage_6[12][3]), .b(stage_6[12][4]), .cin(stage_6[12][5]), .cout(stage_7[13][1]), .s(stage_7[12][3]) );
assign stage_7[12][4] = stage_6[12][6];
FA FA_7_21 ( .a(stage_6[13][0]), .b(stage_6[13][1]), .cin(stage_6[13][2]), .cout(stage_7[14][0]), .s(stage_7[13][2]) );
FA FA_7_22 ( .a(stage_6[13][3]), .b(stage_6[13][4]), .cin(stage_6[13][5]), .cout(stage_7[14][1]), .s(stage_7[13][3]) );
assign stage_7[13][4] = stage_6[13][6];
FA FA_7_23 ( .a(stage_6[14][0]), .b(stage_6[14][1]), .cin(stage_6[14][2]), .cout(stage_7[15][0]), .s(stage_7[14][2]) );
FA FA_7_24 ( .a(stage_6[14][3]), .b(stage_6[14][4]), .cin(stage_6[14][5]), .cout(stage_7[15][1]), .s(stage_7[14][3]) );
assign stage_7[14][4] = stage_6[14][6];
FA FA_7_25 ( .a(stage_6[15][0]), .b(stage_6[15][1]), .cin(stage_6[15][2]), .cout(stage_7[16][0]), .s(stage_7[15][2]) );
FA FA_7_26 ( .a(stage_6[15][3]), .b(stage_6[15][4]), .cin(stage_6[15][5]), .cout(stage_7[16][1]), .s(stage_7[15][3]) );
assign stage_7[15][4] = stage_6[15][6];
FA FA_7_27 ( .a(stage_6[16][0]), .b(stage_6[16][1]), .cin(stage_6[16][2]), .cout(stage_7[17][0]), .s(stage_7[16][2]) );
FA FA_7_28 ( .a(stage_6[16][3]), .b(stage_6[16][4]), .cin(stage_6[16][5]), .cout(stage_7[17][1]), .s(stage_7[16][3]) );
assign stage_7[16][4] = stage_6[16][6];
FA FA_7_29 ( .a(stage_6[17][0]), .b(stage_6[17][1]), .cin(stage_6[17][2]), .cout(stage_7[18][0]), .s(stage_7[17][2]) );
FA FA_7_30 ( .a(stage_6[17][3]), .b(stage_6[17][4]), .cin(stage_6[17][5]), .cout(stage_7[18][1]), .s(stage_7[17][3]) );
FA FA_7_31 ( .a(stage_6[18][0]), .b(stage_6[18][1]), .cin(stage_6[18][2]), .cout(stage_7[19][0]), .s(stage_7[18][2]) );
HA HA_7_2 ( .a(stage_6[18][3]), .b(stage_6[18][4]), .cout(stage_7[19][1]), .s(stage_7[18][3]) );
FA FA_7_32 ( .a(stage_6[19][0]), .b(stage_6[19][1]), .cin(stage_6[19][2]), .cout(stage_7[20][0]), .s(stage_7[19][2]) );
assign stage_7[20][1] = stage_6[20][0];

wire stage_8 [`NBIT+8:0][`NDATA*2:0];
assign stage_8[0][0] = stage_7[0][0];
assign stage_8[1][0] = stage_7[1][0];
FA FA_8_0 ( .a(stage_7[2][0]), .b(stage_7[2][1]), .cin(stage_7[2][2]), .cout(stage_8[3][0]), .s(stage_8[2][0]) );
FA FA_8_1 ( .a(stage_7[3][0]), .b(stage_7[3][1]), .cin(stage_7[3][2]), .cout(stage_8[4][0]), .s(stage_8[3][1]) );
assign stage_8[3][2] = stage_7[3][3];
FA FA_8_2 ( .a(stage_7[4][0]), .b(stage_7[4][1]), .cin(stage_7[4][2]), .cout(stage_8[5][0]), .s(stage_8[4][1]) );
HA HA_8_0 ( .a(stage_7[4][3]), .b(stage_7[4][4]), .cout(stage_8[5][1]), .s(stage_8[4][2]) );
FA FA_8_3 ( .a(stage_7[5][0]), .b(stage_7[5][1]), .cin(stage_7[5][2]), .cout(stage_8[6][0]), .s(stage_8[5][2]) );
FA FA_8_4 ( .a(stage_7[5][3]), .b(stage_7[5][4]), .cin(stage_7[5][5]), .cout(stage_8[6][1]), .s(stage_8[5][3]) );
FA FA_8_5 ( .a(stage_7[6][0]), .b(stage_7[6][1]), .cin(stage_7[6][2]), .cout(stage_8[7][0]), .s(stage_8[6][2]) );
HA HA_8_1 ( .a(stage_7[6][3]), .b(stage_7[6][4]), .cout(stage_8[7][1]), .s(stage_8[6][3]) );
FA FA_8_6 ( .a(stage_7[7][0]), .b(stage_7[7][1]), .cin(stage_7[7][2]), .cout(stage_8[8][0]), .s(stage_8[7][2]) );
HA HA_8_2 ( .a(stage_7[7][3]), .b(stage_7[7][4]), .cout(stage_8[8][1]), .s(stage_8[7][3]) );
FA FA_8_7 ( .a(stage_7[8][0]), .b(stage_7[8][1]), .cin(stage_7[8][2]), .cout(stage_8[9][0]), .s(stage_8[8][2]) );
HA HA_8_3 ( .a(stage_7[8][3]), .b(stage_7[8][4]), .cout(stage_8[9][1]), .s(stage_8[8][3]) );
FA FA_8_8 ( .a(stage_7[9][0]), .b(stage_7[9][1]), .cin(stage_7[9][2]), .cout(stage_8[10][0]), .s(stage_8[9][2]) );
HA HA_8_4 ( .a(stage_7[9][3]), .b(stage_7[9][4]), .cout(stage_8[10][1]), .s(stage_8[9][3]) );
FA FA_8_9 ( .a(stage_7[10][0]), .b(stage_7[10][1]), .cin(stage_7[10][2]), .cout(stage_8[11][0]), .s(stage_8[10][2]) );
HA HA_8_5 ( .a(stage_7[10][3]), .b(stage_7[10][4]), .cout(stage_8[11][1]), .s(stage_8[10][3]) );
FA FA_8_10 ( .a(stage_7[11][0]), .b(stage_7[11][1]), .cin(stage_7[11][2]), .cout(stage_8[12][0]), .s(stage_8[11][2]) );
HA HA_8_6 ( .a(stage_7[11][3]), .b(stage_7[11][4]), .cout(stage_8[12][1]), .s(stage_8[11][3]) );
FA FA_8_11 ( .a(stage_7[12][0]), .b(stage_7[12][1]), .cin(stage_7[12][2]), .cout(stage_8[13][0]), .s(stage_8[12][2]) );
HA HA_8_7 ( .a(stage_7[12][3]), .b(stage_7[12][4]), .cout(stage_8[13][1]), .s(stage_8[12][3]) );
FA FA_8_12 ( .a(stage_7[13][0]), .b(stage_7[13][1]), .cin(stage_7[13][2]), .cout(stage_8[14][0]), .s(stage_8[13][2]) );
HA HA_8_8 ( .a(stage_7[13][3]), .b(stage_7[13][4]), .cout(stage_8[14][1]), .s(stage_8[13][3]) );
FA FA_8_13 ( .a(stage_7[14][0]), .b(stage_7[14][1]), .cin(stage_7[14][2]), .cout(stage_8[15][0]), .s(stage_8[14][2]) );
HA HA_8_9 ( .a(stage_7[14][3]), .b(stage_7[14][4]), .cout(stage_8[15][1]), .s(stage_8[14][3]) );
FA FA_8_14 ( .a(stage_7[15][0]), .b(stage_7[15][1]), .cin(stage_7[15][2]), .cout(stage_8[16][0]), .s(stage_8[15][2]) );
HA HA_8_10 ( .a(stage_7[15][3]), .b(stage_7[15][4]), .cout(stage_8[16][1]), .s(stage_8[15][3]) );
FA FA_8_15 ( .a(stage_7[16][0]), .b(stage_7[16][1]), .cin(stage_7[16][2]), .cout(stage_8[17][0]), .s(stage_8[16][2]) );
HA HA_8_11 ( .a(stage_7[16][3]), .b(stage_7[16][4]), .cout(stage_8[17][1]), .s(stage_8[16][3]) );
FA FA_8_16 ( .a(stage_7[17][0]), .b(stage_7[17][1]), .cin(stage_7[17][2]), .cout(stage_8[18][0]), .s(stage_8[17][2]) );
assign stage_8[17][3] = stage_7[17][3];
FA FA_8_17 ( .a(stage_7[18][0]), .b(stage_7[18][1]), .cin(stage_7[18][2]), .cout(stage_8[19][0]), .s(stage_8[18][1]) );
assign stage_8[18][2] = stage_7[18][3];
FA FA_8_18 ( .a(stage_7[19][0]), .b(stage_7[19][1]), .cin(stage_7[19][2]), .cout(stage_8[20][0]), .s(stage_8[19][1]) );
HA HA_8_12 ( .a(stage_7[20][0]), .b(stage_7[20][1]), .cout(stage_8[21][0]), .s(stage_8[20][1]) );

wire stage_9 [`NBIT+9:0][`NDATA*2:0];
assign stage_9[0][0] = stage_8[0][0];
assign stage_9[1][0] = stage_8[1][0];
assign stage_9[2][0] = stage_8[2][0];
FA FA_9_0 ( .a(stage_8[3][0]), .b(stage_8[3][1]), .cin(stage_8[3][2]), .cout(stage_9[4][0]), .s(stage_9[3][0]) );
FA FA_9_1 ( .a(stage_8[4][0]), .b(stage_8[4][1]), .cin(stage_8[4][2]), .cout(stage_9[5][0]), .s(stage_9[4][1]) );
FA FA_9_2 ( .a(stage_8[5][0]), .b(stage_8[5][1]), .cin(stage_8[5][2]), .cout(stage_9[6][0]), .s(stage_9[5][1]) );
assign stage_9[5][2] = stage_8[5][3];
FA FA_9_3 ( .a(stage_8[6][0]), .b(stage_8[6][1]), .cin(stage_8[6][2]), .cout(stage_9[7][0]), .s(stage_9[6][1]) );
assign stage_9[6][2] = stage_8[6][3];
FA FA_9_4 ( .a(stage_8[7][0]), .b(stage_8[7][1]), .cin(stage_8[7][2]), .cout(stage_9[8][0]), .s(stage_9[7][1]) );
assign stage_9[7][2] = stage_8[7][3];
FA FA_9_5 ( .a(stage_8[8][0]), .b(stage_8[8][1]), .cin(stage_8[8][2]), .cout(stage_9[9][0]), .s(stage_9[8][1]) );
assign stage_9[8][2] = stage_8[8][3];
FA FA_9_6 ( .a(stage_8[9][0]), .b(stage_8[9][1]), .cin(stage_8[9][2]), .cout(stage_9[10][0]), .s(stage_9[9][1]) );
assign stage_9[9][2] = stage_8[9][3];
FA FA_9_7 ( .a(stage_8[10][0]), .b(stage_8[10][1]), .cin(stage_8[10][2]), .cout(stage_9[11][0]), .s(stage_9[10][1]) );
assign stage_9[10][2] = stage_8[10][3];
FA FA_9_8 ( .a(stage_8[11][0]), .b(stage_8[11][1]), .cin(stage_8[11][2]), .cout(stage_9[12][0]), .s(stage_9[11][1]) );
assign stage_9[11][2] = stage_8[11][3];
FA FA_9_9 ( .a(stage_8[12][0]), .b(stage_8[12][1]), .cin(stage_8[12][2]), .cout(stage_9[13][0]), .s(stage_9[12][1]) );
assign stage_9[12][2] = stage_8[12][3];
FA FA_9_10 ( .a(stage_8[13][0]), .b(stage_8[13][1]), .cin(stage_8[13][2]), .cout(stage_9[14][0]), .s(stage_9[13][1]) );
assign stage_9[13][2] = stage_8[13][3];
FA FA_9_11 ( .a(stage_8[14][0]), .b(stage_8[14][1]), .cin(stage_8[14][2]), .cout(stage_9[15][0]), .s(stage_9[14][1]) );
assign stage_9[14][2] = stage_8[14][3];
FA FA_9_12 ( .a(stage_8[15][0]), .b(stage_8[15][1]), .cin(stage_8[15][2]), .cout(stage_9[16][0]), .s(stage_9[15][1]) );
assign stage_9[15][2] = stage_8[15][3];
FA FA_9_13 ( .a(stage_8[16][0]), .b(stage_8[16][1]), .cin(stage_8[16][2]), .cout(stage_9[17][0]), .s(stage_9[16][1]) );
assign stage_9[16][2] = stage_8[16][3];
FA FA_9_14 ( .a(stage_8[17][0]), .b(stage_8[17][1]), .cin(stage_8[17][2]), .cout(stage_9[18][0]), .s(stage_9[17][1]) );
assign stage_9[17][2] = stage_8[17][3];
FA FA_9_15 ( .a(stage_8[18][0]), .b(stage_8[18][1]), .cin(stage_8[18][2]), .cout(stage_9[19][0]), .s(stage_9[18][1]) );
HA HA_9_0 ( .a(stage_8[19][0]), .b(stage_8[19][1]), .cout(stage_9[20][0]), .s(stage_9[19][1]) );
HA HA_9_1 ( .a(stage_8[20][0]), .b(stage_8[20][1]), .cout(stage_9[21][0]), .s(stage_9[20][1]) );

wire stage_10 [`NBIT+10:0][`NDATA*2:0];
assign stage_10[0][0] = stage_9[0][0];
assign stage_10[1][0] = stage_9[1][0];
assign stage_10[2][0] = stage_9[2][0];
assign stage_10[3][0] = stage_9[3][0];
HA HA_10_0 ( .a(stage_9[4][0]), .b(stage_9[4][1]), .cout(stage_10[5][0]), .s(stage_10[4][0]) );
FA FA_10_0 ( .a(stage_9[5][0]), .b(stage_9[5][1]), .cin(stage_9[5][2]), .cout(stage_10[6][0]), .s(stage_10[5][1]) );
FA FA_10_1 ( .a(stage_9[6][0]), .b(stage_9[6][1]), .cin(stage_9[6][2]), .cout(stage_10[7][0]), .s(stage_10[6][1]) );
FA FA_10_2 ( .a(stage_9[7][0]), .b(stage_9[7][1]), .cin(stage_9[7][2]), .cout(stage_10[8][0]), .s(stage_10[7][1]) );
FA FA_10_3 ( .a(stage_9[8][0]), .b(stage_9[8][1]), .cin(stage_9[8][2]), .cout(stage_10[9][0]), .s(stage_10[8][1]) );
FA FA_10_4 ( .a(stage_9[9][0]), .b(stage_9[9][1]), .cin(stage_9[9][2]), .cout(stage_10[10][0]), .s(stage_10[9][1]) );
FA FA_10_5 ( .a(stage_9[10][0]), .b(stage_9[10][1]), .cin(stage_9[10][2]), .cout(stage_10[11][0]), .s(stage_10[10][1]) );
FA FA_10_6 ( .a(stage_9[11][0]), .b(stage_9[11][1]), .cin(stage_9[11][2]), .cout(stage_10[12][0]), .s(stage_10[11][1]) );
FA FA_10_7 ( .a(stage_9[12][0]), .b(stage_9[12][1]), .cin(stage_9[12][2]), .cout(stage_10[13][0]), .s(stage_10[12][1]) );
FA FA_10_8 ( .a(stage_9[13][0]), .b(stage_9[13][1]), .cin(stage_9[13][2]), .cout(stage_10[14][0]), .s(stage_10[13][1]) );
FA FA_10_9 ( .a(stage_9[14][0]), .b(stage_9[14][1]), .cin(stage_9[14][2]), .cout(stage_10[15][0]), .s(stage_10[14][1]) );
FA FA_10_10 ( .a(stage_9[15][0]), .b(stage_9[15][1]), .cin(stage_9[15][2]), .cout(stage_10[16][0]), .s(stage_10[15][1]) );
FA FA_10_11 ( .a(stage_9[16][0]), .b(stage_9[16][1]), .cin(stage_9[16][2]), .cout(stage_10[17][0]), .s(stage_10[16][1]) );
FA FA_10_12 ( .a(stage_9[17][0]), .b(stage_9[17][1]), .cin(stage_9[17][2]), .cout(stage_10[18][0]), .s(stage_10[17][1]) );
HA HA_10_1 ( .a(stage_9[18][0]), .b(stage_9[18][1]), .cout(stage_10[19][0]), .s(stage_10[18][1]) );
HA HA_10_2 ( .a(stage_9[19][0]), .b(stage_9[19][1]), .cout(stage_10[20][0]), .s(stage_10[19][1]) );
HA HA_10_3 ( .a(stage_9[20][0]), .b(stage_9[20][1]), .cout(stage_10[21][0]), .s(stage_10[20][1]) );

wire [20:0] rca_co;
assign o_result[0] = stage_10[0][0];
assign rca_co[0] = 1'b0;
FA FA_final_1( .a(stage_10[1][0]), .b(1'b0), .cin(rca_co[0]), .cout(rca_co[1]), .s(o_result[1]) );
FA FA_final_2( .a(stage_10[2][0]), .b(1'b0), .cin(rca_co[1]), .cout(rca_co[2]), .s(o_result[2]) );
FA FA_final_3( .a(stage_10[3][0]), .b(1'b0), .cin(rca_co[2]), .cout(rca_co[3]), .s(o_result[3]) );
FA FA_final_4( .a(stage_10[4][0]), .b(1'b0), .cin(rca_co[3]), .cout(rca_co[4]), .s(o_result[4]) );
FA FA_final_5( .a(stage_10[5][0]), .b(stage_10[5][1]), .cin(rca_co[4]), .cout(rca_co[5]), .s(o_result[5]) );
FA FA_final_6( .a(stage_10[6][0]), .b(stage_10[6][1]), .cin(rca_co[5]), .cout(rca_co[6]), .s(o_result[6]) );
FA FA_final_7( .a(stage_10[7][0]), .b(stage_10[7][1]), .cin(rca_co[6]), .cout(rca_co[7]), .s(o_result[7]) );
FA FA_final_8( .a(stage_10[8][0]), .b(stage_10[8][1]), .cin(rca_co[7]), .cout(rca_co[8]), .s(o_result[8]) );
FA FA_final_9( .a(stage_10[9][0]), .b(stage_10[9][1]), .cin(rca_co[8]), .cout(rca_co[9]), .s(o_result[9]) );
FA FA_final_10( .a(stage_10[10][0]), .b(stage_10[10][1]), .cin(rca_co[9]), .cout(rca_co[10]), .s(o_result[10]) );
FA FA_final_11( .a(stage_10[11][0]), .b(stage_10[11][1]), .cin(rca_co[10]), .cout(rca_co[11]), .s(o_result[11]) );
FA FA_final_12( .a(stage_10[12][0]), .b(stage_10[12][1]), .cin(rca_co[11]), .cout(rca_co[12]), .s(o_result[12]) );
FA FA_final_13( .a(stage_10[13][0]), .b(stage_10[13][1]), .cin(rca_co[12]), .cout(rca_co[13]), .s(o_result[13]) );
FA FA_final_14( .a(stage_10[14][0]), .b(stage_10[14][1]), .cin(rca_co[13]), .cout(rca_co[14]), .s(o_result[14]) );
FA FA_final_15( .a(stage_10[15][0]), .b(stage_10[15][1]), .cin(rca_co[14]), .cout(rca_co[15]), .s(o_result[15]) );
FA FA_final_16( .a(stage_10[16][0]), .b(stage_10[16][1]), .cin(rca_co[15]), .cout(rca_co[16]), .s(o_result[16]) );
FA FA_final_17( .a(stage_10[17][0]), .b(stage_10[17][1]), .cin(rca_co[16]), .cout(rca_co[17]), .s(o_result[17]) );
FA FA_final_18( .a(stage_10[18][0]), .b(stage_10[18][1]), .cin(rca_co[17]), .cout(rca_co[18]), .s(o_result[18]) );
FA FA_final_19( .a(stage_10[19][0]), .b(stage_10[19][1]), .cin(rca_co[18]), .cout(rca_co[19]), .s(o_result[19]) );
FA FA_final_20( .a(stage_10[20][0]), .b(stage_10[20][1]), .cin(rca_co[19]), .cout(rca_co[20]), .s(o_result[20]) );
FA FA_final_21( .a(stage_10[21][0]), .b(1'b0), .cin(rca_co[20]), .cout(o_result[22]), .s(o_result[21]) );

endmodule